magic
tech tsmc180
timestamp 1701440386
<< nwell >>
rect 0 618 297 1323
<< polysilicon >>
rect 110 780 119 798
rect 148 780 157 798
rect 110 645 119 682
rect 148 646 157 682
rect 110 588 119 624
rect 148 588 157 625
rect 110 523 119 534
rect 148 523 157 534
<< ndiffusion >>
rect 107 534 110 588
rect 119 534 148 588
rect 157 534 160 588
<< pdiffusion >>
rect 107 682 110 780
rect 119 682 123 780
rect 145 682 148 780
rect 157 682 160 780
<< ntransistor >>
rect 110 534 119 588
rect 148 534 157 588
<< ptransistor >>
rect 110 682 119 780
rect 148 682 157 780
<< polycontact >>
rect 104 624 125 645
rect 142 625 163 646
<< ndiffcontact >>
rect 86 534 107 588
rect 160 534 181 588
<< pdiffcontact >>
rect 85 682 107 780
rect 123 682 145 780
rect 160 682 182 780
<< psubstratetap >>
rect 169 16 204 51
<< nsubstratetap >>
rect 117 1285 152 1320
<< metal1 >>
rect 0 1320 297 1323
rect 0 1312 117 1320
rect 0 1293 56 1312
rect 75 1293 117 1312
rect 0 1285 117 1293
rect 152 1311 297 1320
rect 152 1292 190 1311
rect 209 1292 297 1311
rect 152 1285 297 1292
rect 0 1283 297 1285
rect 0 1259 297 1271
rect 0 1232 297 1244
rect 77 1191 107 1213
rect 85 780 107 1191
rect 160 1190 187 1212
rect 160 780 182 1190
rect 129 670 141 682
rect 129 658 187 670
rect 175 639 187 658
rect 175 627 227 639
rect 175 613 187 627
rect 166 601 187 613
rect 166 588 178 601
rect 86 187 107 534
rect 81 166 107 187
rect 0 128 297 140
rect 0 99 297 111
rect 0 70 297 82
rect 0 51 297 54
rect 0 46 169 51
rect 0 27 60 46
rect 79 27 169 46
rect 0 16 169 27
rect 204 16 297 51
rect 0 14 297 16
<< m2contact >>
rect 56 1293 75 1312
rect 190 1292 209 1311
rect 55 1191 77 1213
rect 187 1190 209 1212
rect 104 624 125 645
rect 142 625 163 646
rect 227 624 246 643
rect 60 167 81 186
rect 60 27 79 46
<< metal2 >>
rect 58 1213 72 1293
rect 99 1276 113 1337
rect 132 1304 146 1337
rect 132 1290 160 1304
rect 99 1262 121 1276
rect 107 645 121 1262
rect 146 646 160 1290
rect 192 1212 206 1292
rect 231 643 245 1337
rect 62 46 76 167
rect 107 75 121 624
rect 99 61 121 75
rect 99 0 113 61
rect 146 47 160 625
rect 132 33 160 47
rect 132 0 146 33
rect 231 0 245 624
<< labels >>
rlabel metal1 0 14 0 54 3 GND!
rlabel metal1 0 70 0 82 3 nReset
rlabel metal1 0 99 0 111 3 Clock
rlabel metal1 0 128 0 140 3 Test
rlabel metal1 0 1283 0 1323 3 Vdd!
rlabel metal1 0 1259 0 1271 3 ScanReturn
rlabel metal1 0 1232 0 1244 3 Scan
rlabel metal2 99 1337 113 1337 5 A
rlabel metal2 132 1337 146 1337 5 B
rlabel metal2 231 1337 245 1337 5 Y
rlabel metal2 132 0 146 0 1 B
rlabel metal1 297 1283 297 1323 7 Vdd!
rlabel metal1 297 1259 297 1271 7 ScanReturn
rlabel metal1 297 1232 297 1244 7 Scan
rlabel metal2 231 0 245 0 1 Y
rlabel metal1 297 128 297 140 7 Test
rlabel metal1 297 99 297 111 7 Clock
rlabel metal1 297 70 297 82 7 nReset
rlabel metal1 297 14 297 54 7 GND!
rlabel metal2 99 0 113 0 1 A
<< end >>
