magic
tech tsmc180
timestamp 1701337852
<< nwell >>
rect 0 412 848 1339
<< polysilicon >>
rect 95 734 104 827
rect 166 734 175 822
rect 237 734 246 822
rect 314 734 323 823
rect 386 734 395 823
rect 455 734 464 820
rect 524 734 533 820
rect 670 734 679 820
rect 95 224 104 636
rect 166 529 175 636
rect 166 330 175 431
rect 237 403 246 636
rect 314 529 323 636
rect 166 224 175 276
rect 237 224 246 382
rect 314 370 323 431
rect 386 373 395 636
rect 455 590 464 636
rect 393 352 395 373
rect 314 330 323 349
rect 314 224 323 276
rect 386 224 395 352
rect 455 224 464 569
rect 524 564 533 636
rect 670 618 679 636
rect 677 597 679 618
rect 524 224 533 543
rect 670 257 679 597
rect 670 224 679 236
rect 95 61 104 170
rect 166 147 175 170
rect 166 58 175 126
rect 237 118 246 170
rect 314 118 323 170
rect 386 118 395 170
rect 455 118 464 170
rect 524 154 533 170
rect 670 150 679 170
<< ndiffusion >>
rect 163 276 166 330
rect 175 276 178 330
rect 311 276 314 330
rect 323 276 327 330
rect 92 170 95 224
rect 104 170 166 224
rect 175 170 212 224
rect 233 170 237 224
rect 246 170 314 224
rect 323 170 359 224
rect 380 170 386 224
rect 395 170 398 224
rect 419 170 455 224
rect 464 170 524 224
rect 533 170 536 224
rect 667 170 670 224
rect 679 170 682 224
<< pdiffusion >>
rect 92 636 95 734
rect 104 636 113 734
rect 134 636 166 734
rect 175 636 192 734
rect 213 636 237 734
rect 246 636 254 734
rect 275 636 314 734
rect 323 636 340 734
rect 361 636 386 734
rect 395 636 415 734
rect 436 636 455 734
rect 464 636 484 734
rect 505 636 524 734
rect 533 636 536 734
rect 667 636 670 734
rect 679 636 682 734
rect 163 431 166 529
rect 175 431 178 529
rect 311 431 314 529
rect 323 431 326 529
<< ntransistor >>
rect 166 276 175 330
rect 314 276 323 330
rect 95 170 104 224
rect 166 170 175 224
rect 237 170 246 224
rect 314 170 323 224
rect 386 170 395 224
rect 455 170 464 224
rect 524 170 533 224
rect 670 170 679 224
<< ptransistor >>
rect 95 636 104 734
rect 166 636 175 734
rect 237 636 246 734
rect 314 636 323 734
rect 386 636 395 734
rect 455 636 464 734
rect 524 636 533 734
rect 670 636 679 734
rect 166 431 175 529
rect 314 431 323 529
<< polycontact >>
rect 74 556 95 577
rect 225 382 246 403
rect 443 569 464 590
rect 302 349 323 370
rect 372 352 393 373
rect 656 597 677 618
rect 523 543 544 564
rect 658 236 679 257
rect 154 126 175 147
<< ndiffcontact >>
rect 142 276 163 330
rect 178 276 199 330
rect 290 276 311 330
rect 327 276 348 330
rect 71 170 92 224
rect 212 170 233 224
rect 359 170 380 224
rect 398 170 419 224
rect 536 170 557 224
rect 646 170 667 224
rect 682 170 703 224
<< pdiffcontact >>
rect 71 636 92 734
rect 113 636 134 734
rect 192 636 213 734
rect 254 636 275 734
rect 340 636 361 734
rect 415 636 436 734
rect 484 636 505 734
rect 536 636 557 734
rect 646 636 667 734
rect 682 636 703 734
rect 142 431 163 529
rect 178 431 199 529
rect 290 431 311 529
rect 326 431 347 529
<< psubstratetap >>
rect 252 19 513 55
<< nsubstratetap >>
rect 136 1293 764 1321
<< metal1 >>
rect 0 1321 848 1328
rect 0 1293 136 1321
rect 764 1293 848 1321
rect 0 1284 848 1293
rect 0 1260 214 1272
rect 0 1233 67 1245
rect 260 815 272 1284
rect 324 1260 848 1272
rect 608 1233 848 1245
rect 260 780 272 796
rect 75 770 207 779
rect 75 767 192 770
rect 75 734 87 767
rect 260 768 304 780
rect 195 734 207 751
rect 260 734 272 768
rect 292 655 304 768
rect 421 759 553 771
rect 346 734 358 751
rect 421 734 433 759
rect 541 734 553 759
rect 608 671 620 1233
rect 682 1205 848 1217
rect 649 734 661 794
rect 682 734 694 1205
rect 121 624 133 636
rect 488 624 500 636
rect 121 612 500 624
rect 541 613 553 636
rect 691 622 703 636
rect 541 601 656 613
rect 690 610 703 622
rect 50 560 74 572
rect 47 349 83 361
rect 47 141 59 349
rect 80 224 92 236
rect 114 145 126 581
rect 147 573 443 585
rect 147 529 159 573
rect 544 547 605 559
rect 296 529 308 541
rect 199 477 290 489
rect 143 330 155 431
rect 213 386 225 398
rect 287 354 302 366
rect 335 368 347 431
rect 335 356 372 368
rect 335 330 347 356
rect 199 282 290 326
rect 181 248 193 276
rect 181 236 227 248
rect 215 224 227 236
rect 361 240 658 252
rect 215 158 227 170
rect 267 158 279 234
rect 361 224 373 240
rect 691 224 703 610
rect 557 187 646 199
rect 405 158 417 170
rect 545 158 557 170
rect 0 129 59 141
rect 128 131 154 143
rect 267 146 417 158
rect 722 141 734 382
rect 722 129 848 141
rect 0 100 848 112
rect 0 71 848 83
rect 0 55 848 59
rect 0 42 252 55
rect 0 23 210 42
rect 229 23 252 42
rect 0 19 252 23
rect 513 52 848 55
rect 513 33 545 52
rect 564 33 848 52
rect 513 19 848 33
rect 0 15 848 19
<< m2contact >>
rect 214 1253 233 1272
rect 67 1229 86 1248
rect 305 1253 324 1272
rect 257 796 276 815
rect 192 751 211 770
rect 341 751 360 770
rect 291 636 310 655
rect 643 794 662 813
rect 605 652 624 671
rect 110 581 129 600
rect 31 560 50 579
rect 83 349 102 368
rect 77 236 96 255
rect 293 541 312 560
rect 605 547 624 566
rect 194 383 213 402
rect 268 351 287 370
rect 263 234 282 253
rect 717 382 736 401
rect 109 126 128 145
rect 212 139 231 158
rect 542 139 561 158
rect 210 23 229 42
rect 545 33 564 52
<< metal2 >>
rect 33 579 47 1339
rect 99 1330 113 1339
rect 99 1316 124 1330
rect 33 0 47 560
rect 68 397 82 1229
rect 110 600 124 1316
rect 233 1257 305 1271
rect 276 796 643 810
rect 211 753 341 767
rect 293 560 307 636
rect 607 566 621 652
rect 68 383 194 397
rect 271 384 717 398
rect 271 370 285 384
rect 102 351 268 365
rect 96 237 263 251
rect 110 25 124 126
rect 212 42 226 139
rect 547 52 561 139
rect 99 11 124 25
rect 99 0 113 11
<< labels >>
rlabel metal1 848 15 848 59 7 GND!
rlabel metal1 0 1284 0 1328 3 Vdd!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 848 71 848 83 7 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 848 100 848 112 7 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 848 129 848 141 7 Test
rlabel metal2 33 0 47 0 1 D
rlabel metal2 99 0 113 0 1 Load
rlabel metal1 0 15 0 59 3 GND!
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 848 1260 848 1272 7 ScanReturn
rlabel metal2 33 1339 47 1339 5 D
rlabel metal2 99 1339 113 1339 5 Load
rlabel metal1 848 1284 848 1328 7 Vdd!
rlabel metal1 848 1233 848 1245 7 Q
rlabel metal1 848 1205 848 1217 7 M
rlabel metal1 0 1233 0 1245 3 SDI
<< end >>
