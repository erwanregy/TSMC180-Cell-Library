magic
tech tsmc180
timestamp 1701361821
<< nwell >>
rect 27 1078 135 1328
<< polysilicon >>
rect 90 1183 99 1200
rect 90 1045 99 1085
rect 90 202 99 1024
rect 90 137 99 148
<< ndiffusion >>
rect 87 148 90 202
rect 99 148 102 202
<< pdiffusion >>
rect 87 1085 90 1183
rect 99 1085 102 1183
<< ntransistor >>
rect 90 148 99 202
<< ptransistor >>
rect 90 1085 99 1183
<< polycontact >>
rect 78 1024 99 1045
<< ndiffcontact >>
rect 66 148 87 202
rect 102 148 123 202
<< pdiffcontact >>
rect 65 1085 87 1183
rect 102 1085 123 1183
<< psubstratetap >>
rect 44 18 79 53
<< nsubstratetap >>
rect 44 1286 79 1321
<< metal1 >>
rect 0 1321 87 1324
rect 0 1286 44 1321
rect 79 1286 87 1321
rect 0 1284 87 1286
rect 0 1260 53 1272
rect 0 1233 29 1245
rect 17 1041 29 1233
rect 41 1073 53 1260
rect 65 1183 87 1284
rect 111 1073 123 1085
rect 41 1061 123 1073
rect 17 1029 78 1041
rect 111 202 123 1061
rect 66 55 87 148
rect 0 53 369 55
rect 0 18 44 53
rect 79 18 369 53
rect 0 15 369 18
<< m2contact >>
rect 369 15 409 55
<< metal2 >>
rect 165 55 565 1339
rect 165 15 369 55
rect 409 15 565 55
rect 165 0 565 15
<< labels >>
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal1 0 1260 0 1272 3 nScan
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 0 15 0 55 3 GND!
rlabel metal2 165 1339 565 1339 5 GND!
rlabel metal2 165 0 565 0 1 GND!
<< end >>
