magic
tech tsmc180
timestamp 1701693720
use leftbuf  leftbuf_0
timestamp 1701621919
transform 1 0 0 0 1 0
box 0 0 2574 1339
use inv  inv_0
timestamp 1701646065
transform 1 0 2574 0 1 0
box 0 0 132 1339
use smux2  smux2_0
timestamp 1701647509
transform 1 0 2706 0 1 0
box 0 0 429 1339
use rdtype  rdtype_0
timestamp 1701631232
transform 1 0 3135 0 1 0
box 0 0 429 1339
use buffer  buffer_0
timestamp 1701647406
transform 1 0 3564 0 1 0
box 0 0 132 1339
<< end >>
