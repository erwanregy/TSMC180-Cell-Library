magic
tech tsmc180
timestamp 1701609707
<< nwell >>
rect 0 605 561 1328
<< polysilicon >>
rect 68 927 77 1003
rect 139 927 148 1003
rect 216 927 225 1003
rect 288 927 297 1003
rect 462 927 471 1013
rect 68 722 77 829
rect 68 346 77 624
rect 139 388 148 829
rect 216 612 225 829
rect 288 714 297 829
rect 462 798 471 829
rect 469 777 471 798
rect 296 693 297 714
rect 68 240 77 292
rect 139 240 148 367
rect 216 240 225 591
rect 288 240 297 693
rect 462 273 471 777
rect 462 240 471 252
rect 68 146 77 186
rect 68 80 77 125
rect 139 118 148 186
rect 216 118 225 186
rect 288 118 297 186
rect 462 150 471 186
<< ndiffusion >>
rect 65 292 68 346
rect 77 292 80 346
rect 65 186 68 240
rect 77 186 114 240
rect 135 186 139 240
rect 148 186 216 240
rect 225 186 261 240
rect 282 186 288 240
rect 297 186 300 240
rect 459 186 462 240
rect 471 186 474 240
<< pdiffusion >>
rect 65 829 68 927
rect 77 829 94 927
rect 115 829 139 927
rect 148 829 156 927
rect 177 829 216 927
rect 225 829 242 927
rect 263 829 288 927
rect 297 829 300 927
rect 459 829 462 927
rect 471 829 474 927
rect 65 624 68 722
rect 77 624 80 722
<< ntransistor >>
rect 68 292 77 346
rect 68 186 77 240
rect 139 186 148 240
rect 216 186 225 240
rect 288 186 297 240
rect 462 186 471 240
<< ptransistor >>
rect 68 829 77 927
rect 139 829 148 927
rect 216 829 225 927
rect 288 829 297 927
rect 462 829 471 927
rect 68 624 77 722
<< polycontact >>
rect 448 777 469 798
rect 275 693 296 714
rect 216 591 237 612
rect 128 367 149 388
rect 450 252 471 273
rect 58 125 79 146
<< ndiffcontact >>
rect 44 292 65 346
rect 80 292 101 346
rect 44 186 65 240
rect 114 186 135 240
rect 261 186 282 240
rect 300 186 321 240
rect 438 186 459 240
rect 474 186 495 240
<< pdiffcontact >>
rect 44 829 65 927
rect 94 829 115 927
rect 156 829 177 927
rect 242 829 263 927
rect 300 829 321 927
rect 438 829 459 927
rect 474 829 495 927
rect 44 624 65 722
rect 80 624 101 722
<< psubstratetap >>
rect 154 19 415 55
<< nsubstratetap >>
rect 38 1293 471 1321
<< metal1 >>
rect 0 1321 561 1328
rect 0 1293 38 1321
rect 471 1293 561 1321
rect 0 1284 561 1293
rect 0 1260 116 1272
rect 0 1244 86 1245
rect 0 1233 72 1244
rect 162 987 174 1284
rect 217 1260 561 1272
rect 474 1205 561 1217
rect 162 975 453 987
rect 162 927 174 975
rect 441 927 453 975
rect 474 927 486 1205
rect 48 793 60 829
rect 97 817 109 829
rect 246 817 258 829
rect 97 805 258 817
rect 303 793 315 829
rect 483 815 495 829
rect 482 803 495 815
rect 48 781 448 793
rect 49 752 157 764
rect 49 722 61 752
rect 214 697 275 709
rect 85 609 97 624
rect 49 597 97 609
rect 49 383 61 597
rect 49 371 128 383
rect 49 346 61 371
rect 50 252 194 264
rect 50 240 62 252
rect 182 174 194 252
rect 267 256 450 268
rect 267 240 279 256
rect 483 240 495 803
rect 304 174 316 186
rect 182 162 316 174
rect 0 129 58 141
rect 79 129 561 141
rect 0 100 561 112
rect 0 71 561 83
rect 0 55 561 59
rect 0 52 154 55
rect 0 33 118 52
rect 137 33 154 52
rect 0 19 154 33
rect 415 54 561 55
rect 415 35 440 54
rect 459 35 561 54
rect 415 19 561 35
rect 0 15 561 19
<< m2contact >>
rect 116 1253 135 1272
rect 72 1225 91 1244
rect 198 1253 217 1272
rect 156 844 175 863
rect 157 750 176 769
rect 195 697 214 716
rect 217 592 236 611
rect 82 306 101 325
rect 116 197 135 216
rect 439 195 458 214
rect 118 33 137 52
rect 440 35 459 54
<< metal2 >>
rect 135 1257 198 1271
rect 91 1225 211 1239
rect 158 769 172 844
rect 197 716 211 1225
rect 231 611 245 1339
rect 236 592 245 611
rect 87 305 101 306
rect 87 291 134 305
rect 120 216 134 291
rect 120 52 134 197
rect 231 0 245 592
rect 442 54 456 195
<< labels >>
rlabel metal1 0 1284 0 1328 3 Vdd!
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 SDI
rlabel metal1 0 15 0 59 3 GND!
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 71 0 83 3 nReset
rlabel metal2 231 1339 245 1339 5 D
rlabel metal2 231 0 245 0 1 D
rlabel metal1 561 15 561 59 7 GND!
rlabel metal1 561 71 561 83 7 nReset
rlabel metal1 561 100 561 112 7 Clock
rlabel metal1 561 129 561 141 7 Test
rlabel metal1 561 1205 561 1217 7 M
rlabel metal1 561 1284 561 1328 7 Vdd!
rlabel metal1 561 1260 561 1272 7 ScanReturn
<< end >>
