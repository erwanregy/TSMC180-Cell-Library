magic
tech tsmc180
timestamp 1701622087
use leftbuf  leftbuf_0
timestamp 1701621919
transform 1 0 0 0 1 0
box 0 0 2574 1339
use nand2  nand2_0
timestamp 1701618993
transform 1 0 2574 0 1 0
box 0 0 297 1339
use nand3  nand3_0
timestamp 1701619048
transform 1 0 2871 0 1 0
box 0 0 297 1339
use rightend  rightend_0
timestamp 1701619147
transform 1 0 3168 0 1 0
box 0 0 565 1339
<< end >>
