magic
tech tsmc180
timestamp 1701631232
<< nwell >>
rect 0 605 429 1324
<< polysilicon >>
rect 53 1158 62 1169
rect 53 1024 62 1076
rect 53 343 62 942
rect 91 709 100 1200
rect 129 1158 138 1169
rect 302 1164 311 1175
rect 129 849 138 1076
rect 215 1024 224 1035
rect 262 1024 271 1111
rect 167 849 176 972
rect 215 849 224 942
rect 262 849 271 942
rect 302 882 311 1082
rect 129 709 138 767
rect 167 709 176 767
rect 215 676 224 767
rect 262 709 271 767
rect 91 556 100 627
rect 129 556 138 627
rect 167 556 176 627
rect 215 540 224 655
rect 262 556 271 627
rect 91 491 100 502
rect 129 453 138 502
rect 167 453 176 502
rect 215 453 224 519
rect 262 453 271 502
rect 302 453 311 861
rect 378 849 387 860
rect 340 709 349 828
rect 378 676 387 767
rect 340 590 349 627
rect 378 590 387 655
rect 386 569 387 590
rect 340 556 349 569
rect 378 540 387 569
rect 53 253 62 289
rect 53 117 62 199
rect 129 88 138 399
rect 167 327 176 399
rect 215 343 224 399
rect 262 343 271 399
rect 167 231 176 306
rect 215 278 224 289
rect 262 214 271 289
rect 302 231 311 432
rect 340 411 349 502
rect 378 444 387 519
rect 378 379 387 390
rect 167 166 176 177
rect 302 166 311 177
<< ndiffusion >>
rect 88 502 91 556
rect 100 502 129 556
rect 138 502 167 556
rect 176 502 179 556
rect 259 502 262 556
rect 271 502 274 556
rect 337 502 340 556
rect 349 502 352 556
rect 126 399 129 453
rect 138 399 167 453
rect 176 399 184 453
rect 205 399 215 453
rect 224 399 262 453
rect 271 399 274 453
rect 50 289 53 343
rect 62 289 65 343
rect 50 199 53 253
rect 62 199 65 253
rect 205 289 215 343
rect 224 289 262 343
rect 271 289 274 343
rect 164 177 167 231
rect 176 177 179 231
rect 375 390 378 444
rect 387 390 390 444
rect 299 177 302 231
rect 311 177 314 231
<< pdiffusion >>
rect 50 1076 53 1158
rect 62 1076 65 1158
rect 50 942 53 1024
rect 62 942 65 1024
rect 126 1076 129 1158
rect 138 1076 141 1158
rect 299 1082 302 1164
rect 311 1082 314 1164
rect 206 942 215 1024
rect 224 942 232 1024
rect 253 942 262 1024
rect 271 942 276 1024
rect 126 767 129 849
rect 138 767 141 849
rect 162 767 167 849
rect 176 767 185 849
rect 206 767 215 849
rect 224 767 238 849
rect 259 767 262 849
rect 271 767 276 849
rect 88 627 91 709
rect 100 627 105 709
rect 126 627 129 709
rect 138 627 142 709
rect 163 627 167 709
rect 176 627 179 709
rect 259 627 262 709
rect 271 627 276 709
rect 375 767 378 849
rect 387 767 390 849
rect 337 627 340 709
rect 349 627 352 709
<< pohmic >>
rect 88 24 91 48
rect 114 24 117 48
rect 140 24 143 48
<< nohmic >>
rect 88 1291 91 1315
rect 114 1291 117 1315
rect 140 1291 143 1315
<< ntransistor >>
rect 91 502 100 556
rect 129 502 138 556
rect 167 502 176 556
rect 262 502 271 556
rect 340 502 349 556
rect 129 399 138 453
rect 167 399 176 453
rect 215 399 224 453
rect 262 399 271 453
rect 53 289 62 343
rect 53 199 62 253
rect 215 289 224 343
rect 262 289 271 343
rect 167 177 176 231
rect 378 390 387 444
rect 302 177 311 231
<< ptransistor >>
rect 53 1076 62 1158
rect 53 942 62 1024
rect 129 1076 138 1158
rect 302 1082 311 1164
rect 215 942 224 1024
rect 262 942 271 1024
rect 129 767 138 849
rect 167 767 176 849
rect 215 767 224 849
rect 262 767 271 849
rect 91 627 100 709
rect 129 627 138 709
rect 167 627 176 709
rect 262 627 271 709
rect 378 767 387 849
rect 340 627 349 709
<< polycontact >>
rect 85 1200 106 1221
rect 252 1111 273 1132
rect 159 972 180 993
rect 291 861 312 882
rect 205 655 226 676
rect 205 519 226 540
rect 328 828 349 849
rect 378 655 399 676
rect 329 569 350 590
rect 365 569 386 590
rect 378 519 399 540
rect 300 432 321 453
rect 47 96 68 117
rect 155 306 176 327
rect 328 390 349 411
rect 252 193 273 214
rect 123 67 144 88
<< ndiffcontact >>
rect 67 502 88 556
rect 179 502 200 556
rect 238 502 259 556
rect 274 502 295 556
rect 316 502 337 556
rect 352 502 373 556
rect 105 399 126 453
rect 184 399 205 453
rect 274 399 295 453
rect 29 289 50 343
rect 65 289 86 343
rect 29 199 50 253
rect 65 199 86 253
rect 184 289 205 343
rect 274 289 295 343
rect 143 177 164 231
rect 179 177 200 231
rect 354 390 375 444
rect 390 390 411 444
rect 278 177 299 231
rect 314 177 335 231
<< pdiffcontact >>
rect 29 1076 50 1158
rect 65 1076 86 1158
rect 29 942 50 1024
rect 65 942 86 1024
rect 105 1076 126 1158
rect 141 1076 162 1158
rect 278 1082 299 1164
rect 314 1082 335 1164
rect 185 942 206 1024
rect 232 942 253 1024
rect 276 942 297 1024
rect 105 767 126 849
rect 141 767 162 849
rect 185 767 206 849
rect 238 767 259 849
rect 276 767 297 849
rect 67 627 88 709
rect 105 627 126 709
rect 142 627 163 709
rect 179 627 200 709
rect 238 627 259 709
rect 276 627 297 709
rect 354 767 375 849
rect 390 767 411 849
rect 316 627 337 709
rect 352 627 373 709
<< psubstratetap >>
rect 65 24 88 48
rect 91 24 114 48
rect 117 24 140 48
rect 143 24 166 48
<< nsubstratetap >>
rect 65 1291 88 1315
rect 91 1291 114 1315
rect 117 1291 140 1315
rect 143 1291 166 1315
<< metal1 >>
rect 0 1315 429 1324
rect 0 1303 65 1315
rect 0 1284 17 1303
rect 36 1291 65 1303
rect 88 1291 91 1315
rect 114 1291 117 1315
rect 140 1291 143 1315
rect 166 1291 429 1315
rect 36 1284 429 1291
rect 0 1260 429 1272
rect 0 1233 363 1245
rect 382 1233 429 1245
rect 0 1205 85 1217
rect 106 1205 429 1217
rect 74 1170 153 1182
rect 17 1059 29 1170
rect 74 1158 86 1170
rect 141 1158 153 1170
rect 162 1115 252 1127
rect 273 1111 278 1132
rect 105 1059 117 1076
rect 314 1059 326 1082
rect 17 1047 326 1059
rect 17 744 29 1047
rect 232 1024 244 1047
rect 86 976 159 988
rect 180 972 185 993
rect 194 930 206 942
rect 280 930 292 942
rect 194 918 292 930
rect 150 894 336 906
rect 150 849 162 894
rect 247 861 291 873
rect 247 849 259 861
rect 324 849 336 894
rect 324 828 328 849
rect 349 828 354 849
rect 105 744 117 767
rect 185 744 197 767
rect 276 744 288 767
rect 390 744 402 767
rect 17 732 402 744
rect 67 709 79 732
rect 142 709 154 732
rect 238 709 250 732
rect 316 709 328 732
rect 200 655 205 676
rect 373 655 378 676
rect 114 615 126 627
rect 179 615 191 627
rect 114 603 191 615
rect 285 615 297 627
rect 352 615 364 627
rect 285 603 364 615
rect 328 590 351 591
rect 328 569 329 590
rect 350 569 351 590
rect 328 568 351 569
rect 364 569 365 590
rect 386 569 387 590
rect 364 568 387 569
rect 200 519 205 540
rect 295 522 316 534
rect 373 519 378 540
rect 67 490 79 502
rect 238 490 250 502
rect 17 478 250 490
rect 17 172 29 478
rect 184 453 196 478
rect 295 432 300 453
rect 114 378 126 399
rect 349 390 354 411
rect 390 378 402 390
rect 114 366 402 378
rect 176 306 184 327
rect 74 277 86 289
rect 274 277 286 289
rect 74 265 286 277
rect 86 219 143 231
rect 273 193 278 214
rect 188 165 200 177
rect 314 165 326 177
rect 188 153 326 165
rect 0 129 429 141
rect 0 100 47 112
rect 68 100 429 112
rect 0 71 123 83
rect 144 71 429 83
rect 0 36 17 55
rect 36 48 429 55
rect 36 36 65 48
rect 0 24 65 36
rect 88 24 91 48
rect 114 24 117 48
rect 140 24 143 48
rect 166 24 429 48
rect 0 15 429 24
<< m2contact >>
rect 17 1284 36 1303
rect 363 1229 382 1248
rect 17 1170 36 1189
rect 330 570 349 589
rect 366 570 385 589
rect 17 153 36 172
rect 17 36 36 55
<< metal2 >>
rect 17 1189 31 1284
rect 330 590 344 1339
rect 363 1248 377 1339
rect 330 589 346 590
rect 363 589 377 1229
rect 363 570 366 589
rect 330 569 346 570
rect 17 55 31 153
rect 330 0 344 569
rect 363 0 377 570
<< labels >>
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 1284 0 1324 1 Vdd!
rlabel metal1 0 1233 0 1245 1 Q
rlabel metal1 0 1260 0 1272 1 ScanReturn
rlabel metal1 0 1205 0 1217 1 D
rlabel metal1 429 1284 429 1324 7 Vdd!
rlabel metal1 429 1205 429 1217 7 D
rlabel metal1 429 1260 429 1272 7 ScanReturn
rlabel metal1 429 129 429 141 1 Test
rlabel metal1 429 100 429 112 1 Clock
rlabel metal1 429 71 429 83 1 nReset
rlabel metal1 429 15 429 55 1 GND!
rlabel metal1 429 1233 429 1245 7 Q
rlabel metal2 330 0 344 0 1 nQ
rlabel metal2 330 1339 344 1339 5 nQ
rlabel metal2 363 0 377 0 1 Q
rlabel metal2 363 1339 377 1339 5 Q
<< end >>
