magic
tech tsmc180
timestamp 1701693217
<< nwell >>
rect 0 605 297 1284
<< polysilicon >>
rect 56 835 65 846
rect 104 835 113 846
rect 56 561 65 736
rect 104 596 113 736
rect 167 704 176 846
rect 221 835 230 846
rect 167 593 176 605
rect 221 593 230 736
rect 56 471 65 488
rect 55 450 65 471
rect 56 431 65 450
rect 56 347 65 358
rect 104 347 113 575
rect 166 572 176 593
rect 167 561 176 572
rect 167 347 176 488
rect 221 431 230 572
rect 221 347 230 358
<< ndiffusion >>
rect 53 540 56 561
rect 32 488 56 540
rect 65 509 89 561
rect 65 488 68 509
rect 32 379 56 431
rect 53 358 56 379
rect 65 410 68 431
rect 65 358 89 410
rect 125 509 167 561
rect 146 488 167 509
rect 176 540 179 561
rect 200 540 201 561
rect 176 488 201 540
rect 197 379 221 431
rect 218 358 221 379
rect 230 410 233 431
rect 230 358 254 410
<< pdiffusion >>
rect 32 757 56 835
rect 53 736 56 757
rect 65 757 104 835
rect 65 736 73 757
rect 94 736 104 757
rect 113 814 116 835
rect 113 736 137 814
rect 216 814 221 835
rect 195 736 221 814
rect 230 757 254 835
rect 230 736 233 757
rect 146 683 167 704
rect 125 605 167 683
rect 176 626 200 704
rect 176 605 179 626
<< ntransistor >>
rect 56 488 65 561
rect 56 358 65 431
rect 167 488 176 561
rect 221 358 230 431
<< ptransistor >>
rect 56 736 65 835
rect 104 736 113 835
rect 221 736 230 835
rect 167 605 176 704
<< polycontact >>
rect 92 575 113 596
rect 34 450 55 471
rect 145 572 166 593
rect 209 572 230 593
<< ndiffcontact >>
rect 32 540 53 561
rect 68 488 89 509
rect 32 358 53 379
rect 68 410 89 431
rect 125 488 146 509
rect 179 540 200 561
rect 197 358 218 379
rect 233 410 254 431
<< pdiffcontact >>
rect 32 736 53 757
rect 73 736 94 757
rect 116 814 137 835
rect 195 814 216 835
rect 233 736 254 757
rect 125 683 146 704
rect 179 605 200 626
<< psubstratetap >>
rect 167 17 204 52
<< nsubstratetap >>
rect 174 1286 209 1321
<< metal1 >>
rect 0 1321 297 1324
rect 0 1306 174 1321
rect 0 1285 125 1306
rect 146 1286 174 1306
rect 209 1286 297 1321
rect 146 1285 297 1286
rect 0 1284 297 1285
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 137 814 195 835
rect 232 757 255 758
rect 32 596 53 736
rect 73 704 94 736
rect 232 736 233 757
rect 254 736 255 757
rect 232 735 255 736
rect 124 704 147 705
rect 73 683 125 704
rect 146 683 147 704
rect 124 682 147 683
rect 91 596 114 597
rect 32 575 92 596
rect 113 575 114 596
rect 32 561 53 575
rect 91 574 114 575
rect 144 593 167 594
rect 144 572 145 593
rect 166 572 167 593
rect 144 571 167 572
rect 179 593 200 605
rect 179 572 209 593
rect 179 561 200 572
rect 124 509 147 510
rect 89 488 125 509
rect 146 488 147 509
rect 33 471 56 472
rect 33 450 34 471
rect 55 450 56 471
rect 33 449 56 450
rect 68 431 89 488
rect 124 487 147 488
rect 232 431 255 432
rect 232 410 233 431
rect 254 410 255 431
rect 232 409 255 410
rect 53 358 197 379
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 54 297 55
rect 0 33 125 54
rect 146 52 297 54
rect 146 33 167 52
rect 0 17 167 33
rect 204 17 297 52
rect 0 15 297 17
<< m2contact >>
rect 125 1285 146 1306
rect 233 736 254 757
rect 125 683 146 704
rect 145 572 166 593
rect 125 488 146 509
rect 34 450 55 471
rect 233 410 254 431
rect 125 33 146 54
<< metal2 >>
rect 33 1305 47 1339
rect 33 1284 72 1305
rect 50 471 71 1284
rect 125 704 146 1285
rect 165 1284 179 1339
rect 231 1305 245 1339
rect 231 1284 254 1305
rect 165 605 181 1284
rect 160 593 181 605
rect 166 572 181 593
rect 55 450 71 471
rect 49 449 71 450
rect 50 55 71 449
rect 33 34 71 55
rect 125 54 146 488
rect 160 55 181 572
rect 233 757 254 1284
rect 233 431 254 736
rect 233 55 254 410
rect 33 0 47 34
rect 165 0 179 55
rect 231 34 254 55
rect 231 0 245 34
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal2 33 0 47 0 1 Enable
rlabel metal2 165 0 179 0 1 A
rlabel metal2 231 0 245 0 1 Y
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal2 33 1339 47 1339 5 Enable
rlabel metal2 231 1339 245 1339 5 Y
rlabel metal2 165 1339 179 1339 5 A
<< end >>