magic
tech tsmc180
timestamp 1701619147
<< nwell >>
rect 0 605 149 1324
<< polysilicon >>
rect 90 714 99 731
rect 90 576 99 616
rect 90 503 99 555
rect 90 438 99 449
<< ndiffusion >>
rect 87 449 90 503
rect 99 449 102 503
<< pdiffusion >>
rect 87 616 90 714
rect 99 616 102 714
<< ntransistor >>
rect 90 449 99 503
<< ptransistor >>
rect 90 616 99 714
<< polycontact >>
rect 78 555 99 576
<< ndiffcontact >>
rect 66 449 87 503
rect 102 449 123 503
<< pdiffcontact >>
rect 65 616 87 714
rect 102 616 123 714
<< psubstratetap >>
rect 44 18 79 53
<< nsubstratetap >>
rect 44 1286 79 1321
<< metal1 >>
rect 0 1321 87 1324
rect 0 1286 44 1321
rect 79 1286 87 1321
rect 0 1284 87 1286
rect 0 1260 53 1272
rect 0 1233 29 1245
rect 17 572 29 1233
rect 41 604 53 1260
rect 65 714 87 1284
rect 111 604 123 616
rect 41 592 123 604
rect 17 560 78 572
rect 111 503 123 592
rect 66 55 87 449
rect 0 53 369 55
rect 0 18 44 53
rect 79 18 369 53
rect 0 15 369 18
<< m2contact >>
rect 369 15 405 55
<< metal2 >>
rect 165 55 565 1339
rect 165 15 369 55
rect 405 15 565 55
rect 165 0 565 15
<< labels >>
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal1 0 1260 0 1272 3 nScan
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 0 15 0 55 3 GND!
rlabel metal2 165 1339 565 1339 5 GND!
rlabel metal2 165 0 565 0 1 GND!
<< end >>
