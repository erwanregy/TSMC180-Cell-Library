magic
tech tsmc180
timestamp 1701532255
use leftbuf  leftbuf_0
timestamp 1701531860
transform 1 0 0 0 1 0
box 0 0 2706 1339
use nand2  nand2_0
timestamp 1701529121
transform 1 0 2706 0 1 0
box 0 0 297 1339
use nand3  nand3_0
timestamp 1701532217
transform 1 0 3003 0 1 0
box 0 0 297 1339
use rightend  rightend_0
timestamp 1701532021
transform 1 0 3296 0 1 0
box 4 0 565 1339
<< end >>
