magic
tech tsmc180
timestamp 1701882920
<< nwell >>
rect 0 719 297 1324
<< polysilicon >>
rect 119 817 128 828
rect 119 707 128 719
rect 119 674 128 686
rect 119 609 128 620
<< ndiffusion >>
rect 116 653 119 674
rect 95 620 119 653
rect 128 641 152 674
rect 128 620 131 641
<< pdiffusion >>
rect 115 796 119 817
rect 94 719 119 796
rect 128 740 155 817
rect 128 719 134 740
<< ntransistor >>
rect 119 620 128 674
<< ptransistor >>
rect 119 719 128 817
<< polycontact >>
rect 108 686 129 707
<< ndiffcontact >>
rect 95 653 116 674
rect 131 620 152 641
<< pdiffcontact >>
rect 94 796 115 817
rect 134 719 155 740
<< psubstratetap >>
rect 169 17 204 52
<< nsubstratetap >>
rect 186 1287 221 1322
<< metal1 >>
rect 0 1322 297 1324
rect 0 1305 186 1322
rect 0 1284 94 1305
rect 115 1287 186 1305
rect 221 1287 297 1322
rect 115 1284 297 1287
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 134 707 155 719
rect 129 686 155 707
rect 152 620 241 641
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 52 241 55
rect 0 17 169 52
rect 204 35 241 52
rect 262 35 297 55
rect 204 17 297 35
rect 0 15 297 17
<< m2contact >>
rect 94 1284 115 1305
rect 94 796 115 817
rect 95 653 116 674
rect 241 620 262 641
rect 241 35 262 55
<< metal2 >>
rect 132 1305 146 1339
rect 132 1284 155 1305
rect 94 817 115 1284
rect 135 722 155 1284
rect 134 674 155 722
rect 116 653 155 674
rect 95 598 116 653
rect 95 577 155 598
rect 135 55 155 577
rect 132 34 155 55
rect 241 55 262 620
rect 132 0 146 34
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal2 132 0 146 0 1 Low
rlabel metal2 132 1339 146 1339 5 Low
<< end >>
