magic
tech tsmc180
timestamp 1701882597
<< nwell >>
rect 0 719 297 1324
<< polysilicon >>
rect 56 948 65 959
rect 104 948 113 959
rect 56 589 65 850
rect 104 624 113 850
rect 167 817 176 959
rect 221 948 230 959
rect 56 459 65 535
rect 56 394 65 405
rect 104 394 113 603
rect 167 589 176 719
rect 221 621 230 850
rect 167 394 176 535
rect 221 459 230 600
rect 221 394 230 405
<< ndiffusion >>
rect 53 568 56 589
rect 32 535 56 568
rect 65 556 89 589
rect 65 535 68 556
rect 32 426 56 459
rect 53 405 56 426
rect 65 438 68 459
rect 65 405 89 438
rect 125 556 167 589
rect 146 535 167 556
rect 176 568 179 589
rect 200 568 201 589
rect 176 535 201 568
rect 197 426 221 459
rect 218 405 221 426
rect 230 438 233 459
rect 230 405 254 438
<< pdiffusion >>
rect 32 871 56 948
rect 53 850 56 871
rect 65 871 104 948
rect 65 850 73 871
rect 94 850 104 871
rect 113 927 116 948
rect 113 850 137 927
rect 216 927 221 948
rect 195 850 221 927
rect 230 871 254 948
rect 230 850 233 871
rect 146 796 167 817
rect 125 719 167 796
rect 176 740 200 817
rect 176 719 179 740
<< ntransistor >>
rect 56 535 65 589
rect 56 405 65 459
rect 167 535 176 589
rect 221 405 230 459
<< ptransistor >>
rect 56 850 65 948
rect 104 850 113 948
rect 221 850 230 948
rect 167 719 176 817
<< polycontact >>
rect 92 603 113 624
rect 35 478 56 499
rect 146 600 167 621
rect 209 600 230 621
<< ndiffcontact >>
rect 32 568 53 589
rect 68 535 89 556
rect 32 405 53 426
rect 68 438 89 459
rect 125 535 146 556
rect 179 568 200 589
rect 197 405 218 426
rect 233 438 254 459
<< pdiffcontact >>
rect 32 850 53 871
rect 73 850 94 871
rect 116 927 137 948
rect 195 927 216 948
rect 233 850 254 871
rect 125 796 146 817
rect 179 719 200 740
<< psubstratetap >>
rect 167 17 204 52
<< nsubstratetap >>
rect 174 1286 209 1321
<< metal1 >>
rect 0 1321 297 1324
rect 0 1305 174 1321
rect 0 1284 125 1305
rect 146 1286 174 1305
rect 209 1286 297 1321
rect 146 1284 297 1286
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 137 927 195 948
rect 32 624 53 850
rect 73 817 94 850
rect 73 796 125 817
rect 32 603 92 624
rect 179 621 200 719
rect 32 589 53 603
rect 179 600 209 621
rect 179 589 200 600
rect 89 535 125 556
rect 68 459 89 535
rect 53 405 197 426
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 34 125 55
rect 146 52 297 55
rect 146 34 167 52
rect 0 17 167 34
rect 204 17 297 52
rect 0 15 297 17
<< m2contact >>
rect 125 1284 146 1305
rect 233 850 254 871
rect 125 796 146 817
rect 146 600 167 621
rect 125 535 146 556
rect 35 478 56 499
rect 233 438 254 459
rect 125 34 146 55
<< metal2 >>
rect 33 1305 47 1339
rect 33 1284 72 1305
rect 50 499 71 1284
rect 125 817 146 1284
rect 165 1284 179 1339
rect 231 1305 245 1339
rect 231 1284 254 1305
rect 165 663 181 1284
rect 160 621 181 663
rect 167 600 181 621
rect 56 478 71 499
rect 50 55 71 478
rect 33 34 71 55
rect 125 55 146 535
rect 160 55 181 600
rect 233 871 254 1284
rect 233 459 254 850
rect 233 55 254 438
rect 33 0 47 34
rect 165 0 179 55
rect 231 34 254 55
rect 231 0 245 34
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal2 33 0 47 0 1 Enable
rlabel metal2 165 0 179 0 1 A
rlabel metal2 231 0 245 0 1 Y
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal2 33 1339 47 1339 5 Enable
rlabel metal2 231 1339 245 1339 5 Y
rlabel metal2 165 1339 179 1339 5 A
<< end >>
