magic
tech tsmc180
timestamp 1701880688
<< nwell >>
rect 0 605 297 1324
<< polysilicon >>
rect 110 780 119 798
rect 148 780 157 798
rect 185 780 194 798
rect 110 636 119 682
rect 148 645 157 682
rect 185 647 194 682
rect 110 551 119 615
rect 148 551 157 624
rect 185 551 194 626
rect 110 486 119 497
rect 148 486 157 497
rect 185 486 194 497
<< ndiffusion >>
rect 107 497 110 551
rect 119 497 148 551
rect 157 497 160 551
rect 181 497 185 551
rect 194 497 197 551
<< pdiffusion >>
rect 107 682 110 780
rect 119 682 123 780
rect 145 682 148 780
rect 157 682 160 780
rect 182 682 185 780
rect 194 682 197 780
<< nohmic >>
rect 117 1319 152 1320
rect 117 1285 152 1286
<< ntransistor >>
rect 110 497 119 551
rect 148 497 157 551
rect 185 497 194 551
<< ptransistor >>
rect 110 682 119 780
rect 148 682 157 780
rect 185 682 194 780
<< polycontact >>
rect 104 615 125 636
rect 142 624 163 645
rect 179 626 200 647
<< ndiffcontact >>
rect 86 497 107 551
rect 160 497 181 551
rect 197 497 218 551
<< pdiffcontact >>
rect 85 682 107 780
rect 123 682 145 780
rect 160 682 182 780
rect 197 682 219 780
<< psubstratetap >>
rect 188 16 223 51
<< nsubstratetap >>
rect 117 1286 152 1319
<< metal1 >>
rect 0 1319 297 1324
rect 0 1312 117 1319
rect 0 1293 56 1312
rect 75 1293 117 1312
rect 0 1286 117 1293
rect 152 1312 297 1319
rect 152 1293 190 1312
rect 209 1293 297 1312
rect 152 1286 297 1293
rect 0 1284 297 1286
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 77 1191 107 1213
rect 85 780 107 1191
rect 160 1190 187 1212
rect 160 780 182 1190
rect 129 670 141 682
rect 207 671 219 682
rect 129 658 189 670
rect 207 659 232 671
rect 177 647 189 658
rect 141 645 164 646
rect 103 636 126 637
rect 103 615 104 636
rect 125 615 126 636
rect 141 624 142 645
rect 163 624 164 645
rect 141 623 164 624
rect 177 626 179 647
rect 220 639 232 659
rect 220 627 246 639
rect 103 614 126 615
rect 177 602 189 626
rect 94 590 189 602
rect 94 551 106 590
rect 220 586 232 627
rect 206 574 232 586
rect 206 551 218 574
rect 160 186 181 497
rect 160 166 181 167
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 51 297 55
rect 0 47 188 51
rect 0 28 161 47
rect 180 28 188 47
rect 0 16 188 28
rect 223 16 297 51
rect 0 15 297 16
<< m2contact >>
rect 56 1293 75 1312
rect 190 1293 209 1312
rect 55 1191 77 1213
rect 187 1190 209 1212
rect 104 615 125 636
rect 142 624 163 645
rect 246 624 265 643
rect 160 167 181 186
rect 161 28 180 47
<< metal2 >>
rect 58 1213 72 1293
rect 99 1276 113 1339
rect 132 1304 146 1339
rect 132 1290 160 1304
rect 190 1292 209 1293
rect 99 1262 121 1276
rect 107 636 121 1262
rect 146 645 160 1290
rect 192 1212 206 1292
rect 231 1179 245 1339
rect 231 1164 264 1179
rect 250 643 264 1164
rect 107 263 121 615
rect 99 249 121 263
rect 99 0 113 249
rect 146 227 160 624
rect 248 267 262 624
rect 132 213 160 227
rect 231 253 262 267
rect 132 0 146 213
rect 163 47 177 167
rect 231 0 245 253
<< labels >>
rlabel metal2 132 0 146 0 1 B
rlabel metal2 99 0 113 0 1 A
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal2 99 1339 113 1339 5 A
rlabel metal2 132 1339 146 1339 5 B
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal2 231 0 245 0 1 Y
rlabel metal2 231 1339 245 1339 5 Y
<< end >>
