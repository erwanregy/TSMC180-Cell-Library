magic
tech tsmc180
timestamp 1701961147
<< nwell >>
rect 0 605 429 1324
<< polysilicon >>
rect 53 1162 62 1173
rect 53 1019 62 1064
rect 53 343 62 921
rect 91 725 100 1200
rect 129 1166 138 1177
rect 302 1164 311 1175
rect 129 872 138 1068
rect 215 1019 224 1030
rect 262 1019 271 1106
rect 167 872 176 973
rect 215 872 224 921
rect 262 872 271 921
rect 302 905 311 1066
rect 129 725 138 774
rect 167 725 176 774
rect 215 676 224 774
rect 262 725 271 774
rect 91 556 100 627
rect 129 556 138 627
rect 167 556 176 627
rect 215 540 224 655
rect 262 556 271 627
rect 91 491 100 502
rect 129 453 138 502
rect 167 453 176 502
rect 215 453 224 519
rect 262 453 271 502
rect 302 453 311 884
rect 378 881 387 892
rect 340 725 349 860
rect 378 676 387 783
rect 340 590 349 627
rect 378 590 387 655
rect 386 569 387 590
rect 340 556 349 569
rect 378 540 387 569
rect 53 253 62 289
rect 53 117 62 199
rect 129 88 138 399
rect 167 327 176 399
rect 215 343 224 399
rect 262 343 271 399
rect 167 231 176 306
rect 215 278 224 289
rect 262 214 271 289
rect 302 231 311 432
rect 340 411 349 502
rect 378 444 387 519
rect 378 379 387 390
rect 167 166 176 177
rect 302 166 311 177
<< ndiffusion >>
rect 88 502 91 556
rect 100 502 129 556
rect 138 502 167 556
rect 176 502 179 556
rect 259 502 262 556
rect 271 502 274 556
rect 337 502 340 556
rect 349 502 352 556
rect 126 399 129 453
rect 138 399 167 453
rect 176 399 184 453
rect 205 399 215 453
rect 224 399 262 453
rect 271 399 274 453
rect 50 289 53 343
rect 62 289 65 343
rect 50 199 53 253
rect 62 199 65 253
rect 205 289 215 343
rect 224 289 262 343
rect 271 289 274 343
rect 164 177 167 231
rect 176 177 179 231
rect 375 390 378 444
rect 387 390 390 444
rect 299 177 302 231
rect 311 177 314 231
<< pdiffusion >>
rect 50 1064 53 1162
rect 62 1064 65 1162
rect 50 921 53 1019
rect 62 921 65 1019
rect 126 1068 129 1166
rect 138 1068 141 1166
rect 299 1066 302 1164
rect 311 1066 314 1164
rect 206 921 215 1019
rect 224 921 232 1019
rect 253 921 262 1019
rect 271 921 276 1019
rect 126 774 129 872
rect 138 774 141 872
rect 162 774 167 872
rect 176 774 185 872
rect 206 774 215 872
rect 224 774 238 872
rect 259 774 262 872
rect 271 774 276 872
rect 88 627 91 725
rect 100 627 105 725
rect 126 627 129 725
rect 138 627 142 725
rect 163 627 167 725
rect 176 627 179 725
rect 259 627 262 725
rect 271 627 276 725
rect 375 783 378 881
rect 387 783 390 881
rect 337 627 340 725
rect 349 627 352 725
<< pohmic >>
rect 88 24 91 48
rect 114 24 117 48
rect 140 24 143 48
<< nohmic >>
rect 88 1291 91 1315
rect 114 1291 117 1315
rect 140 1291 143 1315
<< ntransistor >>
rect 91 502 100 556
rect 129 502 138 556
rect 167 502 176 556
rect 262 502 271 556
rect 340 502 349 556
rect 129 399 138 453
rect 167 399 176 453
rect 215 399 224 453
rect 262 399 271 453
rect 53 289 62 343
rect 53 199 62 253
rect 215 289 224 343
rect 262 289 271 343
rect 167 177 176 231
rect 378 390 387 444
rect 302 177 311 231
<< ptransistor >>
rect 53 1064 62 1162
rect 53 921 62 1019
rect 129 1068 138 1166
rect 302 1066 311 1164
rect 215 921 224 1019
rect 262 921 271 1019
rect 129 774 138 872
rect 167 774 176 872
rect 215 774 224 872
rect 262 774 271 872
rect 91 627 100 725
rect 129 627 138 725
rect 167 627 176 725
rect 262 627 271 725
rect 378 783 387 881
rect 340 627 349 725
<< polycontact >>
rect 85 1200 106 1221
rect 252 1106 273 1132
rect 159 973 180 994
rect 291 884 312 905
rect 205 655 226 676
rect 205 519 226 540
rect 328 860 349 881
rect 378 655 399 676
rect 329 569 350 590
rect 365 569 386 590
rect 378 519 399 540
rect 300 432 321 453
rect 47 96 68 117
rect 155 306 176 327
rect 328 390 349 411
rect 252 193 273 214
rect 123 67 144 88
<< ndiffcontact >>
rect 67 502 88 556
rect 179 502 200 556
rect 238 502 259 556
rect 274 502 295 556
rect 316 502 337 556
rect 352 502 373 556
rect 105 399 126 453
rect 184 399 205 453
rect 274 399 295 453
rect 29 289 50 343
rect 65 289 86 343
rect 29 199 50 253
rect 65 199 86 253
rect 184 289 205 343
rect 274 289 295 343
rect 143 177 164 231
rect 179 177 200 231
rect 354 390 375 444
rect 390 390 411 444
rect 278 177 299 231
rect 314 177 335 231
<< pdiffcontact >>
rect 29 1064 50 1162
rect 65 1064 86 1162
rect 29 921 50 1019
rect 65 921 86 1019
rect 105 1068 126 1166
rect 141 1068 162 1166
rect 278 1066 299 1164
rect 314 1066 335 1164
rect 185 921 206 1019
rect 232 921 253 1019
rect 276 921 297 1019
rect 105 774 126 872
rect 141 774 162 872
rect 185 774 206 872
rect 238 774 259 872
rect 276 774 297 872
rect 67 627 88 725
rect 105 627 126 725
rect 142 627 163 725
rect 179 627 200 725
rect 238 627 259 725
rect 276 627 297 725
rect 354 783 375 881
rect 390 783 411 881
rect 316 627 337 725
rect 352 627 373 725
<< psubstratetap >>
rect 65 24 88 48
rect 91 24 114 48
rect 117 24 140 48
rect 143 24 166 48
<< nsubstratetap >>
rect 65 1291 88 1315
rect 91 1291 114 1315
rect 117 1291 140 1315
rect 143 1291 166 1315
<< metal1 >>
rect 0 1315 429 1324
rect 0 1303 65 1315
rect 0 1284 15 1303
rect 34 1291 65 1303
rect 88 1291 91 1315
rect 114 1291 117 1315
rect 140 1291 143 1315
rect 166 1291 429 1315
rect 34 1284 429 1291
rect 0 1260 429 1272
rect 0 1233 363 1245
rect 382 1233 429 1245
rect 0 1205 85 1217
rect 17 1052 29 1172
rect 162 1115 252 1127
rect 273 1106 278 1132
rect 105 1052 126 1068
rect 314 1052 335 1066
rect 17 1040 335 1052
rect 17 762 29 1040
rect 232 1019 253 1040
rect 86 977 159 989
rect 180 973 185 994
rect 247 884 291 896
rect 247 872 259 884
rect 349 860 354 881
rect 105 762 126 774
rect 185 762 206 774
rect 276 762 297 774
rect 390 762 411 783
rect 17 750 411 762
rect 67 725 88 750
rect 142 725 163 750
rect 238 725 259 750
rect 316 725 337 750
rect 200 655 205 676
rect 373 655 378 676
rect 114 615 126 627
rect 179 615 191 627
rect 114 603 191 615
rect 285 615 297 627
rect 352 615 364 627
rect 285 603 364 615
rect 328 590 351 591
rect 328 569 329 590
rect 350 569 351 590
rect 328 568 351 569
rect 364 590 387 591
rect 364 569 365 590
rect 386 569 387 590
rect 364 568 387 569
rect 200 519 205 540
rect 295 522 316 534
rect 373 519 378 540
rect 67 490 79 502
rect 238 490 250 502
rect 17 478 250 490
rect 17 172 29 478
rect 184 453 196 478
rect 295 432 300 453
rect 114 378 126 399
rect 349 390 354 411
rect 390 378 402 390
rect 114 366 402 378
rect 176 306 184 327
rect 74 277 86 289
rect 274 277 286 289
rect 74 265 286 277
rect 86 219 143 231
rect 273 193 278 214
rect 188 165 200 177
rect 314 165 326 177
rect 188 153 326 165
rect 0 129 429 141
rect 0 100 47 112
rect 68 100 429 112
rect 0 71 123 83
rect 144 71 429 83
rect 0 36 17 55
rect 36 48 429 55
rect 36 36 65 48
rect 0 24 65 36
rect 88 24 91 48
rect 114 24 117 48
rect 140 24 143 48
rect 166 24 429 48
rect 0 15 429 24
<< m2contact >>
rect 15 1284 34 1303
rect 363 1229 382 1248
rect 10 1172 29 1191
rect 67 1138 86 1157
rect 141 1138 160 1157
rect 187 921 206 940
rect 276 921 295 940
rect 143 822 162 841
rect 330 570 349 589
rect 366 570 385 589
rect 17 153 36 172
rect 17 36 36 55
<< metal2 >>
rect 15 1191 29 1284
rect 86 1141 141 1155
rect 206 924 276 938
rect 330 839 344 1339
rect 162 825 344 839
rect 330 590 344 825
rect 363 1248 377 1339
rect 330 589 346 590
rect 363 589 377 1229
rect 363 570 366 589
rect 330 569 346 570
rect 17 55 31 153
rect 330 0 344 569
rect 363 0 377 570
<< labels >>
rlabel metal2 363 1339 377 1339 5 Q
rlabel metal2 363 0 377 0 1 Q
rlabel metal2 330 1339 344 1339 5 nQ
rlabel metal2 330 0 344 0 1 nQ
rlabel metal1 429 1233 429 1245 7 Q
rlabel metal1 429 15 429 55 1 GND!
rlabel metal1 429 71 429 83 1 nReset
rlabel metal1 429 100 429 112 1 Clock
rlabel metal1 429 129 429 141 1 Test
rlabel metal1 429 1260 429 1272 7 ScanReturn
rlabel metal1 429 1284 429 1324 7 Vdd!
rlabel metal1 0 1205 0 1217 1 D
rlabel metal1 0 1260 0 1272 1 ScanReturn
rlabel metal1 0 1233 0 1245 1 Q
rlabel metal1 0 1284 0 1324 1 Vdd!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
<< end >>
