magic
tech tsmc180
timestamp 1701964457
<< nwell >>
rect 0 605 858 1324
<< polysilicon >>
rect 482 1162 491 1173
rect 482 1019 491 1064
rect 68 927 77 1003
rect 139 927 148 1003
rect 216 927 225 1003
rect 288 927 297 1003
rect 363 927 372 1013
rect 68 722 77 829
rect 68 346 77 624
rect 139 388 148 829
rect 216 612 225 829
rect 288 714 297 829
rect 363 798 372 829
rect 370 777 372 798
rect 296 693 297 714
rect 68 240 77 292
rect 139 240 148 367
rect 216 240 225 591
rect 288 240 297 693
rect 363 273 372 777
rect 482 343 491 921
rect 520 725 529 1200
rect 558 1166 567 1177
rect 731 1164 740 1175
rect 558 872 567 1068
rect 644 1019 653 1030
rect 691 1019 700 1106
rect 596 872 605 973
rect 644 872 653 921
rect 691 872 700 921
rect 731 905 740 1066
rect 558 725 567 774
rect 596 725 605 774
rect 644 676 653 774
rect 691 725 700 774
rect 520 556 529 627
rect 558 556 567 627
rect 596 556 605 627
rect 644 540 653 655
rect 691 556 700 627
rect 520 491 529 502
rect 558 453 567 502
rect 596 453 605 502
rect 644 453 653 519
rect 691 453 700 502
rect 731 453 740 884
rect 807 881 816 892
rect 769 725 778 860
rect 807 676 816 783
rect 769 590 778 627
rect 807 590 816 655
rect 815 569 816 590
rect 769 556 778 569
rect 807 540 816 569
rect 482 253 491 289
rect 363 240 372 252
rect 558 240 567 399
rect 596 327 605 399
rect 644 343 653 399
rect 691 343 700 399
rect 644 278 653 289
rect 68 146 77 186
rect 68 80 77 125
rect 139 118 148 186
rect 216 118 225 186
rect 288 118 297 186
rect 363 150 372 186
rect 482 117 491 199
rect 691 214 700 289
rect 731 231 740 432
rect 769 411 778 502
rect 807 444 816 519
rect 807 379 816 390
rect 558 88 567 186
rect 731 166 740 177
<< ndiffusion >>
rect 65 292 68 346
rect 77 292 80 346
rect 517 502 520 556
rect 529 502 558 556
rect 567 502 596 556
rect 605 502 608 556
rect 688 502 691 556
rect 700 502 703 556
rect 766 502 769 556
rect 778 502 781 556
rect 555 399 558 453
rect 567 399 596 453
rect 605 399 613 453
rect 634 399 644 453
rect 653 399 691 453
rect 700 399 703 453
rect 479 289 482 343
rect 491 289 494 343
rect 65 186 68 240
rect 77 186 114 240
rect 135 186 139 240
rect 148 186 216 240
rect 225 186 261 240
rect 282 186 288 240
rect 297 186 300 240
rect 360 186 363 240
rect 372 186 375 240
rect 479 199 482 253
rect 491 199 494 253
rect 634 289 644 343
rect 653 289 691 343
rect 700 289 703 343
rect 555 186 558 240
rect 567 186 570 240
rect 804 390 807 444
rect 816 390 819 444
rect 728 177 731 231
rect 740 177 743 231
<< pdiffusion >>
rect 479 1064 482 1162
rect 491 1064 494 1162
rect 65 829 68 927
rect 77 829 94 927
rect 115 829 139 927
rect 148 829 156 927
rect 177 829 216 927
rect 225 829 242 927
rect 263 829 288 927
rect 297 829 300 927
rect 360 829 363 927
rect 372 829 375 927
rect 479 921 482 1019
rect 491 921 494 1019
rect 65 624 68 722
rect 77 624 80 722
rect 555 1068 558 1166
rect 567 1068 570 1166
rect 728 1066 731 1164
rect 740 1066 743 1164
rect 635 921 644 1019
rect 653 921 661 1019
rect 682 921 691 1019
rect 700 921 705 1019
rect 555 774 558 872
rect 567 774 570 872
rect 591 774 596 872
rect 605 774 614 872
rect 635 774 644 872
rect 653 774 667 872
rect 688 774 691 872
rect 700 774 705 872
rect 517 627 520 725
rect 529 627 534 725
rect 555 627 558 725
rect 567 627 571 725
rect 592 627 596 725
rect 605 627 608 725
rect 688 627 691 725
rect 700 627 705 725
rect 804 783 807 881
rect 816 783 819 881
rect 766 627 769 725
rect 778 627 781 725
<< pohmic >>
rect 517 24 520 48
rect 543 24 546 48
rect 569 24 572 48
<< nohmic >>
rect 517 1291 520 1315
rect 543 1291 546 1315
rect 569 1291 572 1315
<< ntransistor >>
rect 68 292 77 346
rect 520 502 529 556
rect 558 502 567 556
rect 596 502 605 556
rect 691 502 700 556
rect 769 502 778 556
rect 558 399 567 453
rect 596 399 605 453
rect 644 399 653 453
rect 691 399 700 453
rect 482 289 491 343
rect 68 186 77 240
rect 139 186 148 240
rect 216 186 225 240
rect 288 186 297 240
rect 363 186 372 240
rect 482 199 491 253
rect 644 289 653 343
rect 691 289 700 343
rect 558 186 567 240
rect 807 390 816 444
rect 731 177 740 231
<< ptransistor >>
rect 482 1064 491 1162
rect 68 829 77 927
rect 139 829 148 927
rect 216 829 225 927
rect 288 829 297 927
rect 363 829 372 927
rect 482 921 491 1019
rect 68 624 77 722
rect 558 1068 567 1166
rect 731 1066 740 1164
rect 644 921 653 1019
rect 691 921 700 1019
rect 558 774 567 872
rect 596 774 605 872
rect 644 774 653 872
rect 691 774 700 872
rect 520 627 529 725
rect 558 627 567 725
rect 596 627 605 725
rect 691 627 700 725
rect 807 783 816 881
rect 769 627 778 725
<< polycontact >>
rect 514 1200 535 1221
rect 349 777 370 798
rect 275 693 296 714
rect 216 591 237 612
rect 128 367 149 388
rect 681 1106 702 1132
rect 588 973 609 994
rect 720 884 741 905
rect 634 655 655 676
rect 634 519 655 540
rect 757 860 778 881
rect 807 655 828 676
rect 758 569 779 590
rect 794 569 815 590
rect 807 519 828 540
rect 729 432 750 453
rect 351 252 372 273
rect 584 306 605 327
rect 58 125 79 146
rect 757 390 778 411
rect 681 193 702 214
rect 476 96 497 117
rect 552 67 573 88
<< ndiffcontact >>
rect 44 292 65 346
rect 80 292 101 346
rect 496 502 517 556
rect 608 502 629 556
rect 667 502 688 556
rect 703 502 724 556
rect 745 502 766 556
rect 781 502 802 556
rect 534 399 555 453
rect 613 399 634 453
rect 703 399 724 453
rect 458 289 479 343
rect 494 289 515 343
rect 44 186 65 240
rect 114 186 135 240
rect 261 186 282 240
rect 300 186 321 240
rect 339 186 360 240
rect 375 186 396 240
rect 458 199 479 253
rect 494 199 515 253
rect 613 289 634 343
rect 703 289 724 343
rect 534 186 555 240
rect 570 186 591 240
rect 783 390 804 444
rect 819 390 840 444
rect 707 177 728 231
rect 743 177 764 231
<< pdiffcontact >>
rect 458 1064 479 1162
rect 494 1064 515 1162
rect 44 829 65 927
rect 94 829 115 927
rect 156 829 177 927
rect 242 829 263 927
rect 300 829 321 927
rect 339 829 360 927
rect 375 829 396 927
rect 458 921 479 1019
rect 494 921 515 1019
rect 44 624 65 722
rect 80 624 101 722
rect 534 1068 555 1166
rect 570 1068 591 1166
rect 707 1066 728 1164
rect 743 1066 764 1164
rect 614 921 635 1019
rect 661 921 682 1019
rect 705 921 726 1019
rect 534 774 555 872
rect 570 774 591 872
rect 614 774 635 872
rect 667 774 688 872
rect 705 774 726 872
rect 496 627 517 725
rect 534 627 555 725
rect 571 627 592 725
rect 608 627 629 725
rect 667 627 688 725
rect 705 627 726 725
rect 783 783 804 881
rect 819 783 840 881
rect 745 627 766 725
rect 781 627 802 725
<< psubstratetap >>
rect 62 30 382 51
rect 494 24 517 48
rect 520 24 543 48
rect 546 24 569 48
rect 572 24 595 48
<< nsubstratetap >>
rect 38 1293 392 1314
rect 494 1291 517 1315
rect 520 1291 543 1315
rect 546 1291 569 1315
rect 572 1291 595 1315
<< metal1 >>
rect 0 1315 858 1324
rect 0 1314 494 1315
rect 0 1293 38 1314
rect 392 1303 494 1314
rect 392 1293 444 1303
rect 0 1284 444 1293
rect 463 1291 494 1303
rect 517 1291 520 1315
rect 543 1291 546 1315
rect 569 1291 572 1315
rect 595 1291 858 1315
rect 463 1284 858 1291
rect 0 1260 116 1272
rect 0 1244 86 1245
rect 0 1233 72 1244
rect 162 987 174 1284
rect 217 1260 858 1272
rect 429 1233 792 1245
rect 811 1233 858 1245
rect 375 1205 514 1217
rect 162 975 354 987
rect 162 927 174 975
rect 342 927 354 975
rect 375 927 387 1205
rect 446 1052 458 1172
rect 591 1115 681 1127
rect 702 1106 707 1132
rect 534 1052 555 1068
rect 743 1052 764 1066
rect 446 1040 764 1052
rect 48 793 60 829
rect 97 817 109 829
rect 246 817 258 829
rect 97 805 258 817
rect 303 793 315 829
rect 384 815 396 829
rect 383 803 396 815
rect 48 781 349 793
rect 49 752 157 764
rect 49 722 61 752
rect 214 697 275 709
rect 85 609 97 624
rect 49 597 97 609
rect 215 612 238 613
rect 49 383 61 597
rect 215 591 216 612
rect 237 591 238 612
rect 215 590 238 591
rect 49 371 128 383
rect 49 346 61 371
rect 50 252 194 264
rect 50 240 62 252
rect 182 174 194 252
rect 267 256 351 268
rect 267 240 279 256
rect 384 240 396 803
rect 446 762 458 1040
rect 661 1019 682 1040
rect 515 977 588 989
rect 609 973 614 994
rect 676 884 720 896
rect 676 872 688 884
rect 778 860 783 881
rect 534 762 555 774
rect 614 762 635 774
rect 705 762 726 774
rect 819 762 840 783
rect 446 750 840 762
rect 496 725 517 750
rect 571 725 592 750
rect 667 725 688 750
rect 745 725 766 750
rect 629 655 634 676
rect 802 655 807 676
rect 543 615 555 627
rect 608 615 620 627
rect 543 603 620 615
rect 714 615 726 627
rect 781 615 793 627
rect 714 603 793 615
rect 757 590 780 591
rect 757 569 758 590
rect 779 569 780 590
rect 757 568 780 569
rect 793 590 816 591
rect 793 569 794 590
rect 815 569 816 590
rect 793 568 816 569
rect 629 519 634 540
rect 724 522 745 534
rect 802 519 807 540
rect 496 490 508 502
rect 667 490 679 502
rect 446 478 679 490
rect 304 174 316 186
rect 182 162 316 174
rect 446 172 458 478
rect 613 453 625 478
rect 724 432 729 453
rect 543 378 555 399
rect 778 390 783 411
rect 819 378 831 390
rect 543 366 831 378
rect 605 306 613 327
rect 503 277 515 289
rect 703 277 715 289
rect 503 265 715 277
rect 515 219 534 231
rect 702 193 707 214
rect 579 165 591 186
rect 743 165 755 177
rect 579 153 755 165
rect 0 129 58 141
rect 79 129 858 141
rect 0 100 476 112
rect 497 100 858 112
rect 0 71 552 83
rect 573 71 858 83
rect 0 54 446 55
rect 0 52 341 54
rect 0 51 118 52
rect 137 51 341 52
rect 360 51 446 54
rect 0 30 62 51
rect 382 36 446 51
rect 465 48 858 55
rect 465 36 494 48
rect 382 30 494 36
rect 0 24 494 30
rect 517 24 520 48
rect 543 24 546 48
rect 569 24 572 48
rect 595 24 858 48
rect 0 15 858 24
<< m2contact >>
rect 444 1284 463 1303
rect 116 1253 135 1272
rect 72 1225 91 1244
rect 198 1253 217 1272
rect 792 1229 811 1248
rect 439 1172 458 1191
rect 496 1138 515 1157
rect 570 1138 589 1157
rect 156 844 175 863
rect 157 750 176 769
rect 195 697 214 716
rect 217 592 236 611
rect 82 306 101 325
rect 116 197 135 216
rect 616 921 635 940
rect 705 921 724 940
rect 572 822 591 841
rect 759 570 778 589
rect 795 570 814 589
rect 340 195 359 214
rect 446 153 465 172
rect 118 51 137 52
rect 341 51 360 54
rect 118 33 137 51
rect 341 35 360 51
rect 446 36 465 55
<< metal2 >>
rect 135 1257 198 1271
rect 91 1225 211 1239
rect 158 769 172 844
rect 197 716 211 1225
rect 231 611 245 1339
rect 444 1191 458 1284
rect 515 1141 570 1155
rect 635 924 705 938
rect 759 839 773 1339
rect 591 825 773 839
rect 236 592 245 611
rect 87 305 101 306
rect 87 291 134 305
rect 120 216 134 291
rect 120 52 134 197
rect 231 0 245 592
rect 759 590 773 825
rect 792 1248 806 1339
rect 759 589 775 590
rect 792 589 806 1229
rect 792 570 795 589
rect 759 569 775 570
rect 343 54 357 195
rect 446 55 460 153
rect 759 0 773 569
rect 792 0 806 570
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 SDI
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 71 0 83 3 nReset
rlabel metal2 231 1339 245 1339 5 D
rlabel metal2 231 0 245 0 1 D
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal2 792 1339 806 1339 5 Q
rlabel metal2 792 0 806 0 1 Q
rlabel metal2 759 1339 773 1339 5 nQ
rlabel metal2 759 0 773 0 1 nQ
rlabel metal1 858 1233 858 1245 7 Q
rlabel metal1 858 15 858 55 1 GND!
rlabel metal1 858 71 858 83 1 nReset
rlabel metal1 858 100 858 112 1 Clock
rlabel metal1 858 129 858 141 1 Test
rlabel metal1 858 1260 858 1272 7 ScanReturn
rlabel metal1 858 1284 858 1324 7 Vdd!
<< end >>
