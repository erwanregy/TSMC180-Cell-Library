magic
tech tsmc180
timestamp 1701437959
<< nwell >>
rect 0 610 297 1339
<< polysilicon >>
rect 110 780 119 798
rect 148 780 157 798
rect 185 780 194 798
rect 110 623 119 682
rect 148 624 157 682
rect 185 624 194 682
rect 110 566 119 602
rect 148 566 157 603
rect 185 566 194 603
rect 110 501 119 512
rect 148 501 157 512
rect 185 501 194 512
<< ndiffusion >>
rect 107 512 110 566
rect 119 512 148 566
rect 157 512 185 566
rect 194 512 197 566
<< pdiffusion >>
rect 107 682 110 780
rect 119 682 123 780
rect 145 682 148 780
rect 157 682 160 780
rect 182 682 185 780
rect 194 682 197 780
<< nohmic >>
rect 117 1285 152 1286
<< ntransistor >>
rect 110 512 119 566
rect 148 512 157 566
rect 185 512 194 566
<< ptransistor >>
rect 110 682 119 780
rect 148 682 157 780
rect 185 682 194 780
<< polycontact >>
rect 104 602 125 623
rect 142 603 163 624
rect 179 603 200 624
<< ndiffcontact >>
rect 86 512 107 566
rect 197 512 218 566
<< pdiffcontact >>
rect 85 682 107 780
rect 123 682 145 780
rect 160 682 182 780
rect 197 682 219 780
<< psubstratetap >>
rect 188 17 223 52
<< nsubstratetap >>
rect 117 1286 152 1320
<< metal1 >>
rect 0 1320 297 1324
rect 0 1312 117 1320
rect 0 1294 56 1312
rect 75 1294 117 1312
rect 0 1286 117 1294
rect 152 1311 297 1320
rect 152 1293 194 1311
rect 213 1293 297 1311
rect 152 1286 297 1293
rect 0 1284 297 1286
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 54 1153 76 1191
rect 54 1131 107 1153
rect 193 1152 215 1190
rect 85 780 107 1131
rect 160 1130 215 1152
rect 160 780 182 1130
rect 129 648 141 682
rect 201 648 213 682
rect 129 636 224 648
rect 212 617 224 636
rect 212 605 241 617
rect 212 590 224 605
rect 201 578 224 590
rect 201 566 213 578
rect 86 480 107 512
rect 59 459 107 480
rect 59 186 80 459
rect 59 167 60 186
rect 79 167 80 186
rect 59 166 80 167
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 52 297 55
rect 0 47 188 52
rect 0 28 60 47
rect 79 28 188 47
rect 0 17 188 28
rect 223 17 297 52
rect 0 15 297 17
<< m2contact >>
rect 56 1294 75 1312
rect 194 1293 213 1311
rect 55 1191 77 1213
rect 193 1190 215 1212
rect 104 602 125 623
rect 142 603 163 624
rect 179 603 200 624
rect 241 602 260 621
rect 60 167 79 186
rect 60 28 79 47
<< metal2 >>
rect 56 1293 75 1294
rect 58 1213 72 1293
rect 99 1177 113 1339
rect 132 1252 146 1339
rect 132 1238 149 1252
rect 99 1163 121 1177
rect 107 623 121 1163
rect 135 1129 149 1238
rect 165 1175 179 1339
rect 194 1292 213 1293
rect 196 1212 210 1292
rect 165 1161 197 1175
rect 135 1109 160 1129
rect 146 624 160 1109
rect 183 624 197 1161
rect 231 669 245 1339
rect 231 655 256 669
rect 242 621 256 655
rect 79 167 81 186
rect 62 47 76 167
rect 107 141 121 602
rect 99 127 121 141
rect 99 0 113 127
rect 146 113 160 603
rect 132 99 160 113
rect 132 0 146 99
rect 183 84 197 603
rect 242 569 256 602
rect 165 70 197 84
rect 231 554 256 569
rect 165 0 179 70
rect 231 0 245 554
<< labels >>
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal2 132 1339 146 1339 5 B
rlabel metal2 165 1339 179 1339 5 C
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal2 99 1339 113 1339 5 A
rlabel metal2 231 1339 245 1339 5 Y
rlabel metal2 231 0 245 0 1 Y
rlabel metal2 165 0 179 0 1 C
rlabel metal2 132 0 146 0 1 B
rlabel metal2 99 0 113 0 1 A
<< end >>
