magic
tech tsmc180
timestamp 1701882768
<< nwell >>
rect 0 719 297 1324
<< polysilicon >>
rect 119 817 128 828
rect 119 708 128 719
rect 119 675 128 687
rect 119 610 128 621
<< ndiffusion >>
rect 116 654 119 675
rect 95 621 119 654
rect 128 642 152 675
rect 128 621 131 642
<< pdiffusion >>
rect 115 796 119 817
rect 94 719 119 796
rect 128 796 134 817
rect 128 719 155 796
<< ntransistor >>
rect 119 621 128 675
<< ptransistor >>
rect 119 719 128 817
<< polycontact >>
rect 108 687 129 708
<< ndiffcontact >>
rect 95 654 116 675
rect 131 621 152 642
<< pdiffcontact >>
rect 94 796 115 817
rect 134 796 155 817
<< psubstratetap >>
rect 169 17 204 52
<< nsubstratetap >>
rect 186 1287 221 1322
<< metal1 >>
rect 0 1322 297 1324
rect 0 1305 186 1322
rect 0 1284 94 1305
rect 115 1287 186 1305
rect 221 1287 297 1322
rect 115 1284 297 1287
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 95 687 108 708
rect 95 675 116 687
rect 152 621 241 642
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 52 241 55
rect 0 17 169 52
rect 204 35 241 52
rect 262 35 297 55
rect 204 17 297 35
rect 0 15 297 17
<< m2contact >>
rect 94 1284 115 1305
rect 94 796 115 817
rect 241 621 262 642
rect 241 35 262 55
<< metal2 >>
rect 132 1305 146 1339
rect 132 1284 155 1305
rect 94 817 115 1284
rect 135 55 155 1284
rect 132 34 155 55
rect 241 55 262 621
rect 132 0 146 34
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal2 132 0 146 0 1 High
rlabel metal2 132 1339 146 1339 5 High
<< end >>
