magic
tech tsmc180
timestamp 1701430251
<< nwell >>
rect 0 490 432 1284
<< polysilicon >>
rect 39 955 48 966
rect 110 955 119 966
rect 166 955 175 966
rect 274 878 283 964
rect 39 843 48 857
rect 110 843 119 857
rect 166 843 175 857
rect 39 731 48 745
rect 110 731 119 745
rect 166 731 175 745
rect 274 731 283 857
rect 367 653 376 964
rect 39 588 48 633
rect 110 588 119 633
rect 166 588 175 633
rect 274 588 283 633
rect 367 588 376 632
rect 39 477 48 490
rect 110 477 119 490
rect 166 477 175 490
rect 39 456 76 477
rect 110 456 132 477
rect 166 456 198 477
rect 39 444 48 456
rect 110 444 119 456
rect 166 444 175 456
rect 274 444 283 490
rect 367 444 376 490
rect 39 344 48 390
rect 110 344 119 390
rect 166 344 175 390
rect 274 344 283 389
rect 367 344 376 389
rect 39 276 48 290
rect 110 276 119 290
rect 166 276 175 290
rect 39 208 48 222
rect 110 208 119 222
rect 166 208 175 222
rect 274 208 283 289
rect 39 55 48 154
rect 110 55 119 154
rect 166 55 175 154
rect 274 55 283 187
rect 367 55 376 323
<< ndiffusion >>
rect 36 390 39 444
rect 48 390 110 444
rect 119 390 166 444
rect 175 411 219 444
rect 175 390 198 411
rect 271 422 274 444
rect 250 389 274 422
rect 283 410 318 444
rect 283 389 297 410
rect 364 422 367 444
rect 343 389 367 422
rect 376 410 417 444
rect 376 389 396 410
rect 36 290 39 344
rect 48 323 76 344
rect 97 323 110 344
rect 48 290 110 323
rect 119 311 166 344
rect 119 290 132 311
rect 153 290 166 311
rect 175 323 198 344
rect 175 290 219 323
rect 271 323 274 344
rect 250 289 274 323
rect 283 323 297 344
rect 283 289 318 323
rect 36 222 39 276
rect 48 222 110 276
rect 119 243 166 276
rect 119 222 132 243
rect 153 222 166 243
rect 175 222 219 276
rect 36 187 39 208
rect 15 154 39 187
rect 48 176 110 208
rect 48 155 51 176
rect 72 155 110 176
rect 48 154 110 155
rect 119 187 132 208
rect 153 187 166 208
rect 119 154 166 187
rect 175 187 198 208
rect 175 154 219 187
<< pdiffusion >>
rect 15 878 39 955
rect 36 857 39 878
rect 48 934 51 955
rect 72 934 110 955
rect 48 857 110 934
rect 119 878 166 955
rect 119 857 132 878
rect 153 857 166 878
rect 175 878 219 955
rect 175 857 198 878
rect 36 745 39 843
rect 48 745 110 843
rect 119 822 132 843
rect 153 822 166 843
rect 119 745 166 822
rect 175 745 219 843
rect 36 633 39 731
rect 48 654 110 731
rect 48 633 76 654
rect 97 633 110 654
rect 119 710 132 731
rect 153 710 166 731
rect 119 633 166 710
rect 175 654 219 731
rect 175 633 198 654
rect 250 654 274 731
rect 271 633 274 654
rect 283 654 318 731
rect 283 633 297 654
rect 36 490 39 588
rect 48 490 110 588
rect 119 490 166 588
rect 175 567 198 588
rect 175 490 219 567
rect 250 511 274 588
rect 271 490 274 511
rect 283 567 297 588
rect 283 490 318 567
rect 343 511 367 588
rect 364 490 367 511
rect 376 567 396 588
rect 376 490 417 567
<< ntransistor >>
rect 39 390 48 444
rect 110 390 119 444
rect 166 390 175 444
rect 274 389 283 444
rect 367 389 376 444
rect 39 290 48 344
rect 110 290 119 344
rect 166 290 175 344
rect 274 289 283 344
rect 39 222 48 276
rect 110 222 119 276
rect 166 222 175 276
rect 39 154 48 208
rect 110 154 119 208
rect 166 154 175 208
<< ptransistor >>
rect 39 857 48 955
rect 110 857 119 955
rect 166 857 175 955
rect 39 745 48 843
rect 110 745 119 843
rect 166 745 175 843
rect 39 633 48 731
rect 110 633 119 731
rect 166 633 175 731
rect 274 633 283 731
rect 39 490 48 588
rect 110 490 119 588
rect 166 490 175 588
rect 274 490 283 588
rect 367 490 376 588
<< polycontact >>
rect 262 857 283 878
rect 355 632 376 653
rect 76 456 97 477
rect 132 456 153 477
rect 198 456 219 477
rect 355 323 376 344
rect 262 187 283 208
<< ndiffcontact >>
rect 15 390 36 444
rect 198 390 219 411
rect 250 422 271 444
rect 297 389 318 410
rect 343 422 364 444
rect 396 389 417 410
rect 15 290 36 344
rect 76 323 97 344
rect 132 290 153 311
rect 198 323 219 344
rect 250 323 271 344
rect 297 323 318 344
rect 15 222 36 276
rect 132 222 153 243
rect 15 187 36 208
rect 51 155 72 176
rect 132 187 153 208
rect 198 187 219 208
<< pdiffcontact >>
rect 15 857 36 878
rect 51 934 72 955
rect 132 857 153 878
rect 198 857 219 878
rect 15 745 36 843
rect 132 822 153 843
rect 15 633 36 731
rect 76 633 97 654
rect 132 710 153 731
rect 198 633 219 654
rect 250 633 271 654
rect 297 633 318 654
rect 15 490 36 588
rect 198 567 219 588
rect 250 490 271 511
rect 297 567 318 588
rect 343 490 364 511
rect 396 567 417 588
<< psubstratetap >>
rect 234 18 269 53
<< nsubstratetap >>
rect 235 1285 270 1320
<< metal1 >>
rect 0 1320 432 1324
rect 0 1305 235 1320
rect 0 1284 15 1305
rect 36 1284 51 1305
rect 72 1285 235 1305
rect 270 1285 432 1320
rect 72 1284 432 1285
rect 0 1260 432 1272
rect 0 1233 432 1245
rect 36 857 132 878
rect 219 857 262 878
rect 198 843 219 857
rect 153 822 219 843
rect 36 710 132 731
rect 97 633 198 654
rect 219 633 250 654
rect 318 633 355 653
rect 297 632 355 633
rect 297 621 318 632
rect 198 600 318 621
rect 198 588 219 600
rect 36 490 250 511
rect 271 490 343 511
rect 36 423 250 444
rect 271 422 343 444
rect 198 377 219 390
rect 198 356 318 377
rect 297 344 318 356
rect 97 323 198 344
rect 219 323 250 344
rect 318 323 355 344
rect 36 290 132 311
rect 153 222 219 243
rect 198 208 219 222
rect 36 188 132 208
rect 219 187 262 208
rect 0 129 432 141
rect 0 100 432 112
rect 0 71 432 83
rect 0 34 15 55
rect 36 34 51 55
rect 72 53 432 55
rect 72 34 234 53
rect 0 18 234 34
rect 269 18 432 53
rect 0 15 432 18
<< m2contact >>
rect 15 1284 36 1305
rect 51 1284 72 1305
rect 51 934 72 955
rect 15 745 36 843
rect 15 633 36 731
rect 15 490 36 588
rect 297 567 318 588
rect 396 567 417 588
rect 76 456 97 477
rect 132 456 153 477
rect 198 456 219 477
rect 15 390 36 444
rect 297 389 318 410
rect 396 389 417 410
rect 15 290 36 344
rect 15 222 36 276
rect 51 155 72 176
rect 15 34 36 55
rect 51 34 72 55
<< metal2 >>
rect 99 1324 113 1339
rect 15 843 36 1284
rect 98 1284 113 1324
rect 51 955 72 1284
rect 92 920 113 1284
rect 15 731 36 745
rect 15 588 36 633
rect 76 899 113 920
rect 132 966 146 1339
rect 198 966 212 1339
rect 297 966 311 1339
rect 396 966 410 1339
rect 76 477 97 899
rect 15 344 36 390
rect 15 276 36 290
rect 15 55 36 222
rect 76 211 97 456
rect 132 477 153 966
rect 76 190 113 211
rect 51 55 72 155
rect 99 0 113 190
rect 132 55 153 456
rect 198 477 219 966
rect 198 55 219 456
rect 297 588 318 966
rect 297 410 318 567
rect 297 55 318 389
rect 396 588 417 966
rect 396 410 417 567
rect 396 55 417 389
rect 132 0 146 55
rect 198 0 212 55
rect 297 0 311 55
rect 396 0 410 55
<< labels >>
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 0 15 0 55 3 GND!
rlabel metal2 99 0 113 0 1 A
rlabel metal2 99 1339 113 1339 5 A
rlabel metal2 132 0 146 0 1 B
rlabel metal2 132 1339 146 1339 5 B
rlabel metal2 198 0 212 0 1 Cin
rlabel metal2 198 1339 212 1339 5 Cin
rlabel metal2 297 0 311 0 1 Cout
rlabel metal2 297 1339 311 1339 5 Cout
rlabel metal2 396 0 410 0 1 S
rlabel metal2 396 1339 410 1339 5 S
rlabel metal1 432 1284 432 1324 7 Vdd!
rlabel metal1 432 1260 432 1272 7 ScanReturn
rlabel metal1 432 1233 432 1245 7 Scan
rlabel metal1 432 71 432 83 7 nReset
rlabel metal1 432 100 432 112 7 Clock
rlabel metal1 432 129 432 141 7 Test
rlabel metal1 432 15 432 55 7 GND!
<< end >>