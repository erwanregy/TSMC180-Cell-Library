magic
tech tsmc180
timestamp 1701698285
<< nwell >>
rect 0 605 858 1324
<< polysilicon >>
rect 482 1158 491 1169
rect 482 1024 491 1076
rect 68 927 77 1003
rect 139 927 148 1003
rect 216 927 225 1003
rect 288 927 297 1003
rect 363 927 372 1013
rect 68 722 77 829
rect 68 346 77 624
rect 139 388 148 829
rect 216 612 225 829
rect 288 714 297 829
rect 363 798 372 829
rect 370 777 372 798
rect 296 693 297 714
rect 68 240 77 292
rect 139 240 148 367
rect 216 240 225 591
rect 288 240 297 693
rect 363 273 372 777
rect 482 343 491 942
rect 520 709 529 1200
rect 558 1158 567 1169
rect 731 1164 740 1175
rect 558 849 567 1076
rect 644 1024 653 1035
rect 691 1024 700 1111
rect 596 849 605 972
rect 644 849 653 942
rect 691 849 700 942
rect 731 882 740 1082
rect 558 709 567 767
rect 596 709 605 767
rect 644 676 653 767
rect 691 709 700 767
rect 520 556 529 627
rect 558 556 567 627
rect 596 556 605 627
rect 644 540 653 655
rect 691 556 700 627
rect 520 491 529 502
rect 558 453 567 502
rect 596 453 605 502
rect 644 453 653 519
rect 691 453 700 502
rect 731 453 740 861
rect 807 849 816 860
rect 769 709 778 828
rect 807 676 816 767
rect 769 590 778 627
rect 807 590 816 655
rect 815 569 816 590
rect 769 556 778 569
rect 807 540 816 569
rect 482 253 491 289
rect 363 240 372 252
rect 68 146 77 186
rect 68 80 77 125
rect 139 118 148 186
rect 216 118 225 186
rect 288 118 297 186
rect 363 150 372 186
rect 482 117 491 199
rect 558 88 567 399
rect 596 327 605 399
rect 644 343 653 399
rect 691 343 700 399
rect 596 231 605 306
rect 644 278 653 289
rect 691 214 700 289
rect 731 231 740 432
rect 769 411 778 502
rect 807 444 816 519
rect 807 379 816 390
rect 596 166 605 177
rect 731 166 740 177
<< ndiffusion >>
rect 65 292 68 346
rect 77 292 80 346
rect 517 502 520 556
rect 529 502 558 556
rect 567 502 596 556
rect 605 502 608 556
rect 688 502 691 556
rect 700 502 703 556
rect 766 502 769 556
rect 778 502 781 556
rect 555 399 558 453
rect 567 399 596 453
rect 605 399 613 453
rect 634 399 644 453
rect 653 399 691 453
rect 700 399 703 453
rect 479 289 482 343
rect 491 289 494 343
rect 65 186 68 240
rect 77 186 114 240
rect 135 186 139 240
rect 148 186 216 240
rect 225 186 261 240
rect 282 186 288 240
rect 297 186 300 240
rect 360 186 363 240
rect 372 186 375 240
rect 479 199 482 253
rect 491 199 494 253
rect 634 289 644 343
rect 653 289 691 343
rect 700 289 703 343
rect 593 177 596 231
rect 605 177 608 231
rect 804 390 807 444
rect 816 390 819 444
rect 728 177 731 231
rect 740 177 743 231
<< pdiffusion >>
rect 479 1076 482 1158
rect 491 1076 494 1158
rect 479 942 482 1024
rect 491 942 494 1024
rect 65 829 68 927
rect 77 829 94 927
rect 115 829 139 927
rect 148 829 156 927
rect 177 829 216 927
rect 225 829 242 927
rect 263 829 288 927
rect 297 829 300 927
rect 360 829 363 927
rect 372 829 375 927
rect 65 624 68 722
rect 77 624 80 722
rect 555 1076 558 1158
rect 567 1076 570 1158
rect 728 1082 731 1164
rect 740 1082 743 1164
rect 635 942 644 1024
rect 653 942 661 1024
rect 682 942 691 1024
rect 700 942 705 1024
rect 555 767 558 849
rect 567 767 570 849
rect 591 767 596 849
rect 605 767 614 849
rect 635 767 644 849
rect 653 767 667 849
rect 688 767 691 849
rect 700 767 705 849
rect 517 627 520 709
rect 529 627 534 709
rect 555 627 558 709
rect 567 627 571 709
rect 592 627 596 709
rect 605 627 608 709
rect 688 627 691 709
rect 700 627 705 709
rect 804 767 807 849
rect 816 767 819 849
rect 766 627 769 709
rect 778 627 781 709
<< ntransistor >>
rect 68 292 77 346
rect 520 502 529 556
rect 558 502 567 556
rect 596 502 605 556
rect 691 502 700 556
rect 769 502 778 556
rect 558 399 567 453
rect 596 399 605 453
rect 644 399 653 453
rect 691 399 700 453
rect 482 289 491 343
rect 68 186 77 240
rect 139 186 148 240
rect 216 186 225 240
rect 288 186 297 240
rect 363 186 372 240
rect 482 199 491 253
rect 644 289 653 343
rect 691 289 700 343
rect 596 177 605 231
rect 807 390 816 444
rect 731 177 740 231
<< ptransistor >>
rect 482 1076 491 1158
rect 482 942 491 1024
rect 68 829 77 927
rect 139 829 148 927
rect 216 829 225 927
rect 288 829 297 927
rect 363 829 372 927
rect 68 624 77 722
rect 558 1076 567 1158
rect 731 1082 740 1164
rect 644 942 653 1024
rect 691 942 700 1024
rect 558 767 567 849
rect 596 767 605 849
rect 644 767 653 849
rect 691 767 700 849
rect 520 627 529 709
rect 558 627 567 709
rect 596 627 605 709
rect 691 627 700 709
rect 807 767 816 849
rect 769 627 778 709
<< polycontact >>
rect 514 1200 535 1221
rect 349 777 370 798
rect 275 693 296 714
rect 216 591 237 612
rect 128 367 149 388
rect 681 1111 702 1132
rect 588 972 609 993
rect 720 861 741 882
rect 634 655 655 676
rect 634 519 655 540
rect 757 828 778 849
rect 807 655 828 676
rect 758 569 779 590
rect 794 569 815 590
rect 807 519 828 540
rect 729 432 750 453
rect 351 252 372 273
rect 58 125 79 146
rect 476 96 497 117
rect 584 306 605 327
rect 757 390 778 411
rect 681 193 702 214
rect 552 67 573 88
<< ndiffcontact >>
rect 44 292 65 346
rect 80 292 101 346
rect 496 502 517 556
rect 608 502 629 556
rect 667 502 688 556
rect 703 502 724 556
rect 745 502 766 556
rect 781 502 802 556
rect 534 399 555 453
rect 613 399 634 453
rect 703 399 724 453
rect 458 289 479 343
rect 494 289 515 343
rect 44 186 65 240
rect 114 186 135 240
rect 261 186 282 240
rect 300 186 321 240
rect 339 186 360 240
rect 375 186 396 240
rect 458 199 479 253
rect 494 199 515 253
rect 613 289 634 343
rect 703 289 724 343
rect 572 177 593 231
rect 608 177 629 231
rect 783 390 804 444
rect 819 390 840 444
rect 707 177 728 231
rect 743 177 764 231
<< pdiffcontact >>
rect 458 1076 479 1158
rect 494 1076 515 1158
rect 458 942 479 1024
rect 494 942 515 1024
rect 44 829 65 927
rect 94 829 115 927
rect 156 829 177 927
rect 242 829 263 927
rect 300 829 321 927
rect 339 829 360 927
rect 375 829 396 927
rect 44 624 65 722
rect 80 624 101 722
rect 534 1076 555 1158
rect 570 1076 591 1158
rect 707 1082 728 1164
rect 743 1082 764 1164
rect 614 942 635 1024
rect 661 942 682 1024
rect 705 942 726 1024
rect 534 767 555 849
rect 570 767 591 849
rect 614 767 635 849
rect 667 767 688 849
rect 705 767 726 849
rect 496 627 517 709
rect 534 627 555 709
rect 571 627 592 709
rect 608 627 629 709
rect 667 627 688 709
rect 705 627 726 709
rect 783 767 804 849
rect 819 767 840 849
rect 745 627 766 709
rect 781 627 802 709
<< psubstratetap >>
rect 62 30 721 51
<< nsubstratetap >>
rect 38 1293 720 1314
<< metal1 >>
rect 0 1314 858 1324
rect 0 1293 38 1314
rect 720 1293 858 1314
rect 0 1284 446 1293
rect 465 1284 858 1293
rect 0 1260 116 1272
rect 0 1244 86 1245
rect 0 1233 72 1244
rect 162 987 174 1284
rect 217 1260 858 1272
rect 429 1233 792 1245
rect 811 1233 858 1245
rect 375 1205 514 1217
rect 162 975 354 987
rect 162 927 174 975
rect 342 927 354 975
rect 375 927 387 1205
rect 503 1170 582 1182
rect 446 1059 458 1170
rect 503 1158 515 1170
rect 570 1158 582 1170
rect 591 1115 681 1127
rect 702 1111 707 1132
rect 534 1059 546 1076
rect 743 1059 755 1082
rect 446 1047 755 1059
rect 48 793 60 829
rect 97 817 109 829
rect 246 817 258 829
rect 97 805 258 817
rect 303 793 315 829
rect 384 815 396 829
rect 383 803 396 815
rect 48 781 349 793
rect 49 752 157 764
rect 49 722 61 752
rect 214 697 275 709
rect 85 609 97 624
rect 49 597 97 609
rect 215 612 238 613
rect 49 383 61 597
rect 215 591 216 612
rect 237 591 238 612
rect 215 590 238 591
rect 49 371 128 383
rect 49 346 61 371
rect 50 252 194 264
rect 50 240 62 252
rect 182 174 194 252
rect 267 256 351 268
rect 267 240 279 256
rect 384 240 396 803
rect 446 744 458 1047
rect 661 1024 673 1047
rect 515 976 588 988
rect 609 972 614 993
rect 623 930 635 942
rect 709 930 721 942
rect 623 918 721 930
rect 579 894 765 906
rect 579 849 591 894
rect 676 861 720 873
rect 676 849 688 861
rect 753 849 765 894
rect 753 828 757 849
rect 778 828 783 849
rect 534 744 546 767
rect 614 744 626 767
rect 705 744 717 767
rect 819 744 831 767
rect 446 732 831 744
rect 496 709 508 732
rect 571 709 583 732
rect 667 709 679 732
rect 745 709 757 732
rect 629 655 634 676
rect 802 655 807 676
rect 543 615 555 627
rect 608 615 620 627
rect 543 603 620 615
rect 714 615 726 627
rect 781 615 793 627
rect 714 603 793 615
rect 757 590 780 591
rect 757 569 758 590
rect 779 569 780 590
rect 757 568 780 569
rect 793 590 816 591
rect 793 569 794 590
rect 815 569 816 590
rect 793 568 816 569
rect 629 519 634 540
rect 724 522 745 534
rect 802 519 807 540
rect 496 490 508 502
rect 667 490 679 502
rect 446 478 679 490
rect 304 174 316 186
rect 182 162 316 174
rect 446 172 458 478
rect 613 453 625 478
rect 724 432 729 453
rect 543 378 555 399
rect 778 390 783 411
rect 819 378 831 390
rect 543 366 831 378
rect 605 306 613 327
rect 503 277 515 289
rect 703 277 715 289
rect 503 265 715 277
rect 515 219 572 231
rect 702 193 707 214
rect 617 165 629 177
rect 743 165 755 177
rect 617 153 755 165
rect 0 129 58 141
rect 79 129 858 141
rect 0 100 476 112
rect 497 100 858 112
rect 0 71 552 83
rect 573 71 858 83
rect 0 54 446 55
rect 0 52 341 54
rect 0 51 118 52
rect 137 51 341 52
rect 360 51 446 54
rect 465 51 858 55
rect 0 30 62 51
rect 721 30 858 51
rect 0 15 858 30
<< m2contact >>
rect 446 1293 465 1303
rect 446 1284 465 1293
rect 116 1253 135 1272
rect 72 1225 91 1244
rect 198 1253 217 1272
rect 792 1229 811 1248
rect 446 1170 465 1189
rect 156 844 175 863
rect 157 750 176 769
rect 195 697 214 716
rect 217 592 236 611
rect 82 306 101 325
rect 116 197 135 216
rect 759 570 778 589
rect 795 570 814 589
rect 340 195 359 214
rect 446 153 465 172
rect 118 51 137 52
rect 341 51 360 54
rect 446 51 465 55
rect 118 33 137 51
rect 341 35 360 51
rect 446 36 465 51
<< metal2 >>
rect 135 1257 198 1271
rect 91 1225 211 1239
rect 158 769 172 844
rect 197 716 211 1225
rect 231 611 245 1339
rect 446 1189 460 1284
rect 236 592 245 611
rect 87 305 101 306
rect 87 291 134 305
rect 120 216 134 291
rect 120 52 134 197
rect 231 0 245 592
rect 759 590 773 1339
rect 792 1248 806 1339
rect 759 589 775 590
rect 792 589 806 1229
rect 792 570 795 589
rect 759 569 775 570
rect 343 54 357 195
rect 446 55 460 153
rect 759 0 773 569
rect 792 0 806 570
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 SDI
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 71 0 83 3 nReset
rlabel metal2 231 1339 245 1339 5 D
rlabel metal2 231 0 245 0 1 D
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal1 858 1284 858 1324 7 Vdd!
rlabel metal1 858 1260 858 1272 7 ScanReturn
rlabel metal1 858 129 858 141 1 Test
rlabel metal1 858 100 858 112 1 Clock
rlabel metal1 858 71 858 83 1 nReset
rlabel metal1 858 15 858 55 1 GND!
rlabel metal1 858 1233 858 1245 7 Q
rlabel metal2 759 1339 773 1339 5 nQ
rlabel metal2 792 1339 806 1339 5 Q
rlabel metal2 759 0 773 0 1 nQ
rlabel metal2 792 0 806 0 1 Q
<< end >>
