magic
tech tsmc180
timestamp 1701532021
<< nwell >>
rect 4 1074 153 1324
<< polysilicon >>
rect 94 1183 103 1200
rect 94 1045 103 1085
rect 94 202 103 1024
rect 94 137 103 148
<< ndiffusion >>
rect 91 148 94 202
rect 103 148 106 202
<< pdiffusion >>
rect 91 1085 94 1183
rect 103 1085 106 1183
<< ntransistor >>
rect 94 148 103 202
<< ptransistor >>
rect 94 1085 103 1183
<< polycontact >>
rect 82 1024 103 1045
<< ndiffcontact >>
rect 70 148 91 202
rect 106 148 127 202
<< pdiffcontact >>
rect 69 1085 91 1183
rect 106 1085 127 1183
<< psubstratetap >>
rect 48 18 83 53
<< nsubstratetap >>
rect 48 1286 83 1321
<< metal1 >>
rect 4 1321 91 1324
rect 4 1286 48 1321
rect 83 1286 91 1321
rect 4 1284 91 1286
rect 4 1260 57 1272
rect 4 1233 33 1245
rect 21 1041 33 1233
rect 45 1073 57 1260
rect 69 1183 91 1284
rect 115 1073 127 1085
rect 45 1061 127 1073
rect 21 1029 82 1041
rect 115 202 127 1061
rect 70 55 91 148
rect 4 53 369 55
rect 4 18 48 53
rect 83 18 369 53
rect 4 15 369 18
<< m2contact >>
rect 369 15 409 55
<< metal2 >>
rect 165 55 565 1339
rect 165 15 369 55
rect 409 15 565 55
rect 165 0 565 15
<< labels >>
rlabel metal2 165 1339 565 1339 5 GND!
rlabel metal2 165 0 565 0 1 GND!
rlabel metal1 4 1284 4 1324 3 Vdd!
rlabel metal1 4 1260 4 1272 3 nScan
rlabel metal1 4 1233 4 1245 3 Scan
rlabel metal1 4 15 4 55 3 GND!
<< end >>
