magic
tech tsmc180
timestamp 1701965097
<< nwell >>
rect 0 605 297 1324
<< polysilicon >>
rect 56 834 65 845
rect 104 834 113 845
rect 56 475 65 736
rect 104 510 113 736
rect 167 703 176 845
rect 221 834 230 845
rect 167 508 176 605
rect 56 387 65 421
rect 55 362 65 387
rect 56 345 65 362
rect 56 280 65 291
rect 104 280 113 489
rect 166 485 176 508
rect 221 507 230 736
rect 167 475 176 485
rect 167 280 176 421
rect 221 345 230 486
rect 221 280 230 291
<< ndiffusion >>
rect 53 454 56 475
rect 32 421 56 454
rect 65 442 89 475
rect 65 421 68 442
rect 32 312 56 345
rect 53 291 56 312
rect 65 324 68 345
rect 65 291 89 324
rect 125 442 167 475
rect 146 421 167 442
rect 176 454 179 475
rect 200 454 201 475
rect 176 421 201 454
rect 197 312 221 345
rect 218 291 221 312
rect 230 324 233 345
rect 230 291 254 324
<< pdiffusion >>
rect 32 757 56 834
rect 53 736 56 757
rect 65 757 104 834
rect 65 736 73 757
rect 94 736 104 757
rect 113 813 116 834
rect 113 736 137 813
rect 216 813 221 834
rect 195 736 221 813
rect 230 757 254 834
rect 230 736 233 757
rect 146 682 167 703
rect 125 605 167 682
rect 176 626 200 703
rect 176 605 179 626
<< ntransistor >>
rect 56 421 65 475
rect 56 291 65 345
rect 167 421 176 475
rect 221 291 230 345
<< ptransistor >>
rect 56 736 65 834
rect 104 736 113 834
rect 221 736 230 834
rect 167 605 176 703
<< polycontact >>
rect 92 489 113 510
rect 34 364 55 385
rect 145 486 166 507
rect 209 486 230 507
<< ndiffcontact >>
rect 32 454 53 475
rect 68 421 89 442
rect 32 291 53 312
rect 68 324 89 345
rect 125 421 146 442
rect 179 454 200 475
rect 197 291 218 312
rect 233 324 254 345
<< pdiffcontact >>
rect 32 736 53 757
rect 73 736 94 757
rect 116 813 137 834
rect 195 813 216 834
rect 233 736 254 757
rect 125 682 146 703
rect 179 605 200 626
<< psubstratetap >>
rect 167 17 204 52
<< nsubstratetap >>
rect 174 1286 209 1321
<< metal1 >>
rect 0 1321 297 1324
rect 0 1305 174 1321
rect 0 1284 125 1305
rect 146 1286 174 1305
rect 209 1286 297 1321
rect 146 1284 297 1286
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 137 813 195 834
rect 232 757 255 758
rect 32 510 53 736
rect 73 703 94 736
rect 232 736 233 757
rect 254 736 255 757
rect 232 735 255 736
rect 124 703 147 704
rect 73 682 125 703
rect 146 682 147 703
rect 124 681 147 682
rect 32 489 92 510
rect 144 507 167 508
rect 32 475 53 489
rect 144 486 145 507
rect 166 486 167 507
rect 144 485 167 486
rect 179 507 200 605
rect 179 486 209 507
rect 179 475 200 486
rect 124 442 147 443
rect 89 421 125 442
rect 146 421 147 442
rect 33 385 56 386
rect 33 364 34 385
rect 55 364 56 385
rect 33 363 56 364
rect 68 345 89 421
rect 124 420 147 421
rect 232 345 255 346
rect 232 324 233 345
rect 254 324 255 345
rect 232 323 255 324
rect 53 291 197 312
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 34 125 55
rect 146 52 297 55
rect 146 34 167 52
rect 0 17 167 34
rect 204 17 297 52
rect 0 15 297 17
<< m2contact >>
rect 125 1284 146 1305
rect 233 736 254 757
rect 125 682 146 703
rect 145 486 166 507
rect 125 421 146 442
rect 34 364 55 385
rect 233 324 254 345
rect 125 34 146 55
<< metal2 >>
rect 33 1305 47 1339
rect 33 1284 72 1305
rect 50 387 71 1284
rect 125 703 146 1284
rect 165 1284 179 1339
rect 231 1305 245 1339
rect 231 1284 254 1305
rect 165 549 181 1284
rect 160 508 181 549
rect 159 507 181 508
rect 166 486 181 507
rect 159 485 181 486
rect 49 385 71 387
rect 55 364 71 385
rect 49 362 71 364
rect 50 55 71 362
rect 33 34 71 55
rect 125 55 146 421
rect 160 55 181 485
rect 233 757 254 1284
rect 233 345 254 736
rect 233 55 254 324
rect 33 0 47 34
rect 165 0 179 55
rect 231 34 254 55
rect 231 0 245 34
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal2 33 0 47 0 1 Enable
rlabel metal2 165 0 179 0 1 A
rlabel metal2 231 0 245 0 1 Y
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal2 33 1339 47 1339 5 Enable
rlabel metal2 231 1339 245 1339 5 Y
rlabel metal2 165 1339 179 1339 5 A
<< end >>
