magic
tech tsmc180
timestamp 1701441008
<< nwell >>
rect 0 633 297 1284
<< polysilicon >>
rect 56 863 65 874
rect 104 863 113 874
rect 56 589 65 764
rect 104 624 113 764
rect 167 732 176 874
rect 221 863 230 874
rect 56 459 65 516
rect 56 375 65 386
rect 104 375 113 603
rect 167 589 176 633
rect 221 621 230 764
rect 167 375 176 516
rect 221 459 230 600
rect 221 375 230 386
<< ndiffusion >>
rect 53 568 56 589
rect 32 516 56 568
rect 65 537 89 589
rect 65 516 68 537
rect 32 407 56 459
rect 53 386 56 407
rect 65 438 68 459
rect 65 386 89 438
rect 125 537 167 589
rect 146 516 167 537
rect 176 568 179 589
rect 200 568 201 589
rect 176 516 201 568
rect 197 407 221 459
rect 218 386 221 407
rect 230 438 233 459
rect 230 386 254 438
<< pdiffusion >>
rect 32 785 56 863
rect 53 764 56 785
rect 65 785 104 863
rect 65 764 73 785
rect 94 764 104 785
rect 113 842 116 863
rect 113 764 137 842
rect 216 842 221 863
rect 195 764 221 842
rect 230 785 254 863
rect 230 764 233 785
rect 146 711 167 732
rect 125 633 167 711
rect 176 654 200 732
rect 176 633 179 654
<< ntransistor >>
rect 56 516 65 589
rect 56 386 65 459
rect 167 516 176 589
rect 221 386 230 459
<< ptransistor >>
rect 56 764 65 863
rect 104 764 113 863
rect 221 764 230 863
rect 167 633 176 732
<< polycontact >>
rect 92 603 113 624
rect 35 478 56 499
rect 146 600 167 621
rect 209 600 230 621
<< ndiffcontact >>
rect 32 568 53 589
rect 68 516 89 537
rect 32 386 53 407
rect 68 438 89 459
rect 125 516 146 537
rect 179 568 200 589
rect 197 386 218 407
rect 233 438 254 459
<< pdiffcontact >>
rect 32 764 53 785
rect 73 764 94 785
rect 116 842 137 863
rect 195 842 216 863
rect 233 764 254 785
rect 125 711 146 732
rect 179 633 200 654
<< psubstratetap >>
rect 167 17 204 52
<< nsubstratetap >>
rect 174 1286 209 1321
<< metal1 >>
rect 0 1321 297 1324
rect 0 1305 174 1321
rect 0 1284 125 1305
rect 146 1286 174 1305
rect 209 1286 297 1321
rect 146 1284 297 1286
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 137 842 195 863
rect 32 624 53 764
rect 73 732 94 764
rect 73 711 125 732
rect 32 603 92 624
rect 179 621 200 633
rect 32 589 53 603
rect 179 600 209 621
rect 179 589 200 600
rect 89 516 125 537
rect 68 459 89 516
rect 53 386 197 407
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 34 125 55
rect 146 52 297 55
rect 146 34 167 52
rect 0 17 167 34
rect 204 17 297 52
rect 0 15 297 17
<< m2contact >>
rect 125 1284 146 1305
rect 233 764 254 785
rect 125 711 146 732
rect 146 600 167 621
rect 125 516 146 537
rect 35 478 56 499
rect 233 438 254 459
rect 125 34 146 55
<< metal2 >>
rect 33 1305 47 1339
rect 33 1284 72 1305
rect 50 499 71 1284
rect 125 732 146 1284
rect 165 1284 179 1339
rect 231 1305 245 1339
rect 231 1284 254 1305
rect 165 633 181 1284
rect 160 621 181 633
rect 167 600 181 621
rect 56 478 71 499
rect 50 55 71 478
rect 33 34 71 55
rect 125 55 146 516
rect 160 55 181 600
rect 233 785 254 1284
rect 233 459 254 764
rect 233 55 254 438
rect 33 0 47 34
rect 165 0 179 55
rect 231 34 254 55
rect 231 0 245 34
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal2 33 0 47 0 1 Enable
rlabel metal2 165 0 179 0 1 A
rlabel metal2 231 0 245 0 1 Y
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal2 33 1339 47 1339 5 Enable
rlabel metal2 231 1339 245 1339 5 Y
rlabel metal2 165 1339 179 1339 5 A
<< end >>