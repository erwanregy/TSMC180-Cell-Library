magic
tech tsmc180
timestamp 1701540732
<< nwell >>
rect 0 605 429 1324
<< polysilicon >>
rect 53 1158 62 1169
rect 53 1024 62 1076
rect 53 343 62 942
rect 91 709 100 1200
rect 129 1158 138 1169
rect 302 1164 311 1175
rect 129 849 138 1076
rect 215 1024 224 1035
rect 262 1024 271 1111
rect 167 849 176 972
rect 215 849 224 942
rect 262 849 271 942
rect 302 882 311 1082
rect 129 709 138 767
rect 167 709 176 767
rect 215 676 224 767
rect 262 709 271 767
rect 91 558 100 627
rect 129 558 138 627
rect 167 558 176 627
rect 215 542 224 655
rect 262 558 271 627
rect 91 493 100 504
rect 129 454 138 504
rect 167 454 176 504
rect 215 454 224 521
rect 262 454 271 504
rect 302 454 311 861
rect 378 849 387 860
rect 340 709 349 828
rect 378 676 387 767
rect 340 591 349 627
rect 378 591 387 655
rect 386 570 387 591
rect 340 558 349 570
rect 378 542 387 570
rect 53 253 62 289
rect 53 117 62 199
rect 129 88 138 400
rect 167 327 176 400
rect 215 343 224 400
rect 262 343 271 400
rect 167 231 176 306
rect 215 278 224 289
rect 262 214 271 289
rect 302 231 311 433
rect 340 413 349 504
rect 378 446 387 521
rect 378 381 387 392
rect 167 166 176 177
rect 302 166 311 177
<< ndiffusion >>
rect 88 504 91 558
rect 100 504 129 558
rect 138 504 167 558
rect 176 504 179 558
rect 259 504 262 558
rect 271 504 274 558
rect 337 504 340 558
rect 349 504 352 558
rect 126 400 129 454
rect 138 400 167 454
rect 176 400 184 454
rect 205 400 215 454
rect 224 400 262 454
rect 271 400 274 454
rect 50 289 53 343
rect 62 289 65 343
rect 50 199 53 253
rect 62 199 65 253
rect 205 289 215 343
rect 224 289 262 343
rect 271 289 274 343
rect 164 177 167 231
rect 176 177 179 231
rect 375 392 378 446
rect 387 392 390 446
rect 299 177 302 231
rect 311 177 314 231
<< pdiffusion >>
rect 50 1076 53 1158
rect 62 1076 65 1158
rect 50 942 53 1024
rect 62 942 65 1024
rect 126 1076 129 1158
rect 138 1076 141 1158
rect 299 1082 302 1164
rect 311 1082 314 1164
rect 206 942 215 1024
rect 224 942 232 1024
rect 253 942 262 1024
rect 271 942 276 1024
rect 126 767 129 849
rect 138 767 141 849
rect 162 767 167 849
rect 176 767 185 849
rect 206 767 215 849
rect 224 767 238 849
rect 259 767 262 849
rect 271 767 276 849
rect 88 627 91 709
rect 100 627 105 709
rect 126 627 129 709
rect 138 627 142 709
rect 163 627 167 709
rect 176 627 179 709
rect 259 627 262 709
rect 271 627 276 709
rect 375 767 378 849
rect 387 767 390 849
rect 337 627 340 709
rect 349 627 352 709
<< pohmic >>
rect 88 24 91 48
rect 114 24 117 48
rect 140 24 143 48
<< nohmic >>
rect 88 1291 91 1315
rect 114 1291 117 1315
rect 140 1291 143 1315
<< ntransistor >>
rect 91 504 100 558
rect 129 504 138 558
rect 167 504 176 558
rect 262 504 271 558
rect 340 504 349 558
rect 129 400 138 454
rect 167 400 176 454
rect 215 400 224 454
rect 262 400 271 454
rect 53 289 62 343
rect 53 199 62 253
rect 215 289 224 343
rect 262 289 271 343
rect 167 177 176 231
rect 378 392 387 446
rect 302 177 311 231
<< ptransistor >>
rect 53 1076 62 1158
rect 53 942 62 1024
rect 129 1076 138 1158
rect 302 1082 311 1164
rect 215 942 224 1024
rect 262 942 271 1024
rect 129 767 138 849
rect 167 767 176 849
rect 215 767 224 849
rect 262 767 271 849
rect 91 627 100 709
rect 129 627 138 709
rect 167 627 176 709
rect 262 627 271 709
rect 378 767 387 849
rect 340 627 349 709
<< polycontact >>
rect 85 1200 106 1221
rect 252 1111 273 1132
rect 159 972 180 993
rect 291 861 312 882
rect 205 655 226 676
rect 205 521 226 542
rect 328 828 349 849
rect 378 655 399 676
rect 329 570 350 591
rect 365 570 386 591
rect 378 521 399 542
rect 300 433 321 454
rect 47 96 68 117
rect 155 306 176 327
rect 328 392 349 413
rect 252 193 273 214
rect 123 67 144 88
<< ndiffcontact >>
rect 67 504 88 558
rect 179 504 200 558
rect 238 504 259 558
rect 274 504 295 558
rect 316 504 337 558
rect 352 504 373 558
rect 105 400 126 454
rect 184 400 205 454
rect 274 400 295 454
rect 29 289 50 343
rect 65 289 86 343
rect 29 199 50 253
rect 65 199 86 253
rect 184 289 205 343
rect 274 289 295 343
rect 143 177 164 231
rect 179 177 200 231
rect 354 392 375 446
rect 390 392 411 446
rect 278 177 299 231
rect 314 177 335 231
<< pdiffcontact >>
rect 29 1076 50 1158
rect 65 1076 86 1158
rect 29 942 50 1024
rect 65 942 86 1024
rect 105 1076 126 1158
rect 141 1076 162 1158
rect 278 1082 299 1164
rect 314 1082 335 1164
rect 185 942 206 1024
rect 232 942 253 1024
rect 276 942 297 1024
rect 105 767 126 849
rect 141 767 162 849
rect 185 767 206 849
rect 238 767 259 849
rect 276 767 297 849
rect 67 627 88 709
rect 105 627 126 709
rect 142 627 163 709
rect 179 627 200 709
rect 238 627 259 709
rect 276 627 297 709
rect 354 767 375 849
rect 390 767 411 849
rect 316 627 337 709
rect 352 627 373 709
<< psubstratetap >>
rect 65 24 88 48
rect 91 24 114 48
rect 117 24 140 48
rect 143 24 166 48
<< nsubstratetap >>
rect 65 1291 88 1315
rect 91 1291 114 1315
rect 117 1291 140 1315
rect 143 1291 166 1315
<< metal1 >>
rect 0 1315 429 1324
rect 0 1303 65 1315
rect 0 1284 17 1303
rect 36 1291 65 1303
rect 88 1291 91 1315
rect 114 1291 117 1315
rect 140 1291 143 1315
rect 166 1291 429 1315
rect 36 1284 429 1291
rect 0 1260 429 1272
rect 0 1233 363 1245
rect 382 1233 429 1245
rect 0 1205 85 1217
rect 106 1205 429 1217
rect 74 1170 153 1182
rect 17 1059 29 1170
rect 74 1158 86 1170
rect 141 1158 153 1170
rect 162 1115 252 1127
rect 273 1111 278 1132
rect 105 1059 117 1076
rect 314 1059 326 1082
rect 17 1047 326 1059
rect 17 744 29 1047
rect 232 1024 244 1047
rect 86 976 159 988
rect 180 972 185 993
rect 194 930 206 942
rect 280 930 292 942
rect 194 918 292 930
rect 150 894 336 906
rect 150 849 162 894
rect 247 861 291 873
rect 247 849 259 861
rect 324 849 336 894
rect 324 828 328 849
rect 349 828 354 849
rect 105 744 117 767
rect 185 744 197 767
rect 276 744 288 767
rect 390 744 402 767
rect 17 732 402 744
rect 67 709 79 732
rect 142 709 154 732
rect 238 709 250 732
rect 316 709 328 732
rect 200 655 205 676
rect 373 655 378 676
rect 114 615 126 627
rect 179 615 191 627
rect 114 603 191 615
rect 285 615 297 627
rect 352 615 364 627
rect 285 603 364 615
rect 200 521 205 542
rect 295 524 316 536
rect 373 521 378 542
rect 67 492 79 504
rect 238 492 250 504
rect 17 480 250 492
rect 17 172 29 480
rect 184 454 196 480
rect 295 433 300 454
rect 114 380 126 400
rect 349 392 354 413
rect 390 380 402 392
rect 114 368 402 380
rect 176 306 184 327
rect 74 277 86 289
rect 274 277 286 289
rect 74 265 286 277
rect 86 219 143 231
rect 273 193 278 214
rect 188 165 200 177
rect 314 165 326 177
rect 188 153 326 165
rect 0 129 429 141
rect 0 100 47 112
rect 68 100 429 112
rect 0 71 123 83
rect 144 71 429 83
rect 0 36 17 55
rect 36 48 429 55
rect 36 36 65 48
rect 0 24 65 36
rect 88 24 91 48
rect 114 24 117 48
rect 140 24 143 48
rect 166 24 429 48
rect 0 15 429 24
<< m2contact >>
rect 17 1284 36 1303
rect 363 1229 382 1248
rect 17 1170 36 1189
rect 330 571 349 590
rect 366 571 385 590
rect 17 153 36 172
rect 17 36 36 55
<< metal2 >>
rect 17 1189 31 1284
rect 330 591 344 1339
rect 363 1248 377 1339
rect 330 590 346 591
rect 363 590 377 1229
rect 363 571 366 590
rect 330 570 346 571
rect 17 55 31 153
rect 330 0 344 570
rect 363 0 377 571
<< labels >>
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 1284 0 1324 1 Vdd!
rlabel metal1 0 1233 0 1245 1 Q
rlabel metal1 0 1260 0 1272 1 ScanReturn
rlabel metal1 0 1205 0 1217 1 D
rlabel metal1 429 1284 429 1324 7 Vdd!
rlabel metal1 429 1205 429 1217 7 D
rlabel metal1 429 1260 429 1272 7 ScanReturn
rlabel metal1 429 129 429 141 1 Test
rlabel metal1 429 100 429 112 1 Clock
rlabel metal1 429 71 429 83 1 nReset
rlabel metal1 429 15 429 55 1 GND!
rlabel metal1 429 1233 429 1245 7 Q
rlabel metal2 330 0 344 0 1 nQ
rlabel metal2 330 1339 344 1339 5 nQ
rlabel metal2 363 0 377 0 1 Q
rlabel metal2 363 1339 377 1339 5 Q
<< end >>
