magic
tech tsmc180
timestamp 1701883273
<< nwell >>
rect 0 719 429 1324
<< polysilicon >>
rect 39 1184 48 1195
rect 110 1184 119 1195
rect 166 1184 175 1195
rect 274 1107 283 1193
rect 39 1072 48 1086
rect 110 1072 119 1086
rect 166 1072 175 1086
rect 39 960 48 974
rect 110 960 119 974
rect 166 960 175 974
rect 274 960 283 1086
rect 367 882 376 1193
rect 39 817 48 862
rect 110 817 119 862
rect 166 817 175 862
rect 274 817 283 862
rect 367 817 376 861
rect 39 695 48 719
rect 110 695 119 719
rect 166 695 175 719
rect 39 674 76 695
rect 110 674 132 695
rect 166 674 198 695
rect 39 662 48 674
rect 110 662 119 674
rect 166 662 175 674
rect 274 662 283 719
rect 367 662 376 719
rect 39 562 48 608
rect 110 562 119 608
rect 166 562 175 608
rect 274 562 283 608
rect 367 562 376 608
rect 39 494 48 508
rect 110 494 119 508
rect 166 494 175 508
rect 39 426 48 440
rect 110 426 119 440
rect 166 426 175 440
rect 274 426 283 508
rect 39 55 48 372
rect 110 55 119 372
rect 166 55 175 372
rect 274 55 283 405
rect 367 55 376 541
<< ndiffusion >>
rect 36 608 39 662
rect 48 608 110 662
rect 119 608 166 662
rect 175 629 219 662
rect 175 608 198 629
rect 271 640 274 662
rect 250 608 274 640
rect 283 629 318 662
rect 283 608 297 629
rect 364 640 367 662
rect 343 608 367 640
rect 376 629 417 662
rect 376 608 396 629
rect 36 508 39 562
rect 48 541 76 562
rect 97 541 110 562
rect 48 508 110 541
rect 119 529 166 562
rect 119 508 132 529
rect 153 508 166 529
rect 175 541 198 562
rect 175 508 219 541
rect 271 541 274 562
rect 250 508 274 541
rect 283 541 297 562
rect 283 508 318 541
rect 36 440 39 494
rect 48 440 110 494
rect 119 461 166 494
rect 119 440 132 461
rect 153 440 166 461
rect 175 440 219 494
rect 36 405 39 426
rect 15 372 39 405
rect 48 394 110 426
rect 48 373 51 394
rect 72 373 110 394
rect 48 372 110 373
rect 119 405 132 426
rect 153 405 166 426
rect 119 372 166 405
rect 175 405 198 426
rect 175 372 219 405
<< pdiffusion >>
rect 15 1107 39 1184
rect 36 1086 39 1107
rect 48 1163 51 1184
rect 72 1163 110 1184
rect 48 1086 110 1163
rect 119 1107 166 1184
rect 119 1086 132 1107
rect 153 1086 166 1107
rect 175 1107 219 1184
rect 175 1086 198 1107
rect 36 974 39 1072
rect 48 974 110 1072
rect 119 1051 132 1072
rect 153 1051 166 1072
rect 119 974 166 1051
rect 175 974 219 1072
rect 36 862 39 960
rect 48 883 110 960
rect 48 862 76 883
rect 97 862 110 883
rect 119 939 132 960
rect 153 939 166 960
rect 119 862 166 939
rect 175 883 219 960
rect 175 862 198 883
rect 250 883 274 960
rect 271 862 274 883
rect 283 883 318 960
rect 283 862 297 883
rect 36 719 39 817
rect 48 719 110 817
rect 119 719 166 817
rect 175 796 198 817
rect 175 719 219 796
rect 250 740 274 817
rect 271 719 274 740
rect 283 796 297 817
rect 283 719 318 796
rect 343 740 367 817
rect 364 719 367 740
rect 376 796 396 817
rect 376 719 417 796
<< ntransistor >>
rect 39 608 48 662
rect 110 608 119 662
rect 166 608 175 662
rect 274 608 283 662
rect 367 608 376 662
rect 39 508 48 562
rect 110 508 119 562
rect 166 508 175 562
rect 274 508 283 562
rect 39 440 48 494
rect 110 440 119 494
rect 166 440 175 494
rect 39 372 48 426
rect 110 372 119 426
rect 166 372 175 426
<< ptransistor >>
rect 39 1086 48 1184
rect 110 1086 119 1184
rect 166 1086 175 1184
rect 39 974 48 1072
rect 110 974 119 1072
rect 166 974 175 1072
rect 39 862 48 960
rect 110 862 119 960
rect 166 862 175 960
rect 274 862 283 960
rect 39 719 48 817
rect 110 719 119 817
rect 166 719 175 817
rect 274 719 283 817
rect 367 719 376 817
<< polycontact >>
rect 262 1086 283 1107
rect 355 861 376 882
rect 76 674 97 695
rect 132 674 153 695
rect 198 674 219 695
rect 355 541 376 562
rect 262 405 283 426
<< ndiffcontact >>
rect 15 608 36 662
rect 198 608 219 629
rect 250 640 271 662
rect 297 608 318 629
rect 343 640 364 662
rect 396 608 417 629
rect 15 508 36 562
rect 76 541 97 562
rect 132 508 153 529
rect 198 541 219 562
rect 250 541 271 562
rect 297 541 318 562
rect 15 440 36 494
rect 132 440 153 461
rect 15 405 36 426
rect 51 373 72 394
rect 132 405 153 426
rect 198 405 219 426
<< pdiffcontact >>
rect 15 1086 36 1107
rect 51 1163 72 1184
rect 132 1086 153 1107
rect 198 1086 219 1107
rect 15 974 36 1072
rect 132 1051 153 1072
rect 15 862 36 960
rect 76 862 97 883
rect 132 939 153 960
rect 198 862 219 883
rect 250 862 271 883
rect 297 862 318 883
rect 15 719 36 817
rect 198 796 219 817
rect 250 719 271 740
rect 297 796 318 817
rect 343 719 364 740
rect 396 796 417 817
<< psubstratetap >>
rect 234 18 269 53
<< nsubstratetap >>
rect 235 1285 270 1320
<< metal1 >>
rect 0 1320 429 1324
rect 0 1305 235 1320
rect 0 1284 15 1305
rect 36 1284 51 1305
rect 72 1285 235 1305
rect 270 1285 429 1320
rect 72 1284 429 1285
rect 0 1260 429 1272
rect 0 1233 429 1245
rect 36 1086 132 1107
rect 219 1086 262 1107
rect 198 1072 219 1086
rect 153 1051 219 1072
rect 36 939 132 960
rect 97 862 198 883
rect 219 862 250 883
rect 318 862 355 882
rect 297 861 355 862
rect 297 850 318 861
rect 198 829 318 850
rect 198 817 219 829
rect 36 719 250 740
rect 271 719 343 740
rect 36 641 250 662
rect 271 641 343 662
rect 198 595 219 608
rect 198 574 318 595
rect 297 562 318 574
rect 97 541 198 562
rect 219 541 250 562
rect 318 541 355 562
rect 36 508 132 529
rect 153 440 219 461
rect 198 426 219 440
rect 36 406 132 426
rect 219 405 262 426
rect 0 129 429 141
rect 0 100 429 112
rect 0 71 429 83
rect 0 34 15 55
rect 36 34 51 55
rect 72 53 429 55
rect 72 34 234 53
rect 0 18 234 34
rect 269 18 429 53
rect 0 15 429 18
<< m2contact >>
rect 15 1284 36 1305
rect 51 1284 72 1305
rect 51 1163 72 1184
rect 15 974 36 1072
rect 15 862 36 960
rect 15 719 36 817
rect 297 796 318 817
rect 396 796 417 817
rect 76 674 97 695
rect 132 674 153 695
rect 198 674 219 695
rect 15 608 36 662
rect 297 608 318 629
rect 396 608 417 629
rect 15 508 36 562
rect 15 440 36 494
rect 51 373 72 394
rect 15 34 36 55
rect 51 34 72 55
<< metal2 >>
rect 99 1324 113 1339
rect 15 1072 36 1284
rect 98 1284 113 1324
rect 51 1184 72 1284
rect 92 1149 113 1284
rect 15 960 36 974
rect 15 817 36 862
rect 76 1128 113 1149
rect 132 1195 146 1339
rect 198 1195 212 1339
rect 297 1195 311 1339
rect 396 1195 410 1339
rect 76 695 97 1128
rect 15 562 36 608
rect 15 494 36 508
rect 15 55 36 440
rect 76 429 97 674
rect 132 695 153 1195
rect 76 408 113 429
rect 51 55 72 373
rect 99 0 113 408
rect 132 55 153 674
rect 198 695 219 1195
rect 198 55 219 674
rect 297 817 318 1195
rect 297 629 318 796
rect 297 55 318 608
rect 396 817 417 1195
rect 396 629 417 796
rect 396 55 417 608
rect 132 0 146 55
rect 198 0 212 55
rect 297 0 311 55
rect 396 0 410 55
<< labels >>
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 0 15 0 55 3 GND!
rlabel metal2 99 0 113 0 1 A
rlabel metal2 99 1339 113 1339 5 A
rlabel metal2 132 0 146 0 1 B
rlabel metal2 132 1339 146 1339 5 B
rlabel metal2 198 0 212 0 1 Cin
rlabel metal2 198 1339 212 1339 5 Cin
rlabel metal2 297 0 311 0 1 Cout
rlabel metal2 297 1339 311 1339 5 Cout
rlabel metal2 396 0 410 0 1 S
rlabel metal2 396 1339 410 1339 5 S
rlabel metal1 429 15 429 55 7 GND!
rlabel metal1 429 129 429 141 7 Test
rlabel metal1 429 100 429 112 7 Clock
rlabel metal1 429 71 429 83 7 nReset
rlabel metal1 429 1233 429 1245 7 Scan
rlabel metal1 429 1260 429 1272 7 ScanReturn
rlabel metal1 429 1284 429 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
<< end >>
