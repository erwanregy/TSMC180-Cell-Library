magic
tech tsmc180
timestamp 1701692771
<< nwell >>
rect 0 605 297 1284
<< polysilicon >>
rect 119 706 128 717
rect 119 596 128 607
rect 119 563 128 575
rect 119 498 128 509
<< ndiffusion >>
rect 116 542 119 563
rect 95 509 119 542
rect 128 530 152 563
rect 128 509 131 530
<< pdiffusion >>
rect 115 685 119 706
rect 94 607 119 685
rect 128 685 134 706
rect 128 607 155 685
<< ntransistor >>
rect 119 509 128 563
<< ptransistor >>
rect 119 607 128 706
<< polycontact >>
rect 108 575 129 596
<< ndiffcontact >>
rect 95 542 116 563
rect 131 509 152 530
<< pdiffcontact >>
rect 94 685 115 706
rect 134 685 155 706
<< psubstratetap >>
rect 169 17 204 52
<< nsubstratetap >>
rect 186 1287 221 1322
<< metal1 >>
rect 0 1322 297 1324
rect 0 1306 186 1322
rect 0 1285 94 1306
rect 115 1287 186 1306
rect 221 1287 297 1322
rect 115 1285 297 1287
rect 0 1284 297 1285
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 93 706 116 707
rect 93 685 94 706
rect 115 685 116 706
rect 93 684 116 685
rect 133 706 156 707
rect 133 685 134 706
rect 155 685 156 706
rect 133 684 156 685
rect 95 575 108 596
rect 95 563 116 575
rect 240 530 263 531
rect 152 509 241 530
rect 262 509 263 530
rect 240 508 263 509
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 54 297 55
rect 0 52 241 54
rect 0 17 169 52
rect 204 34 241 52
rect 262 34 297 54
rect 204 17 297 34
rect 0 15 297 17
<< m2contact >>
rect 94 1285 115 1306
rect 94 685 115 706
rect 134 685 155 706
rect 241 509 262 530
rect 241 34 262 54
<< metal2 >>
rect 94 706 115 1285
rect 132 1305 146 1339
rect 132 1284 155 1305
rect 135 706 155 1284
rect 135 55 155 685
rect 132 34 155 55
rect 241 54 262 509
rect 132 0 146 34
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal2 132 0 146 0 1 High
rlabel metal2 132 1339 146 1339 5 High
<< end >>