magic
tech tsmc180
timestamp 1701696883
<< nwell >>
rect 0 605 1056 1324
<< polysilicon >>
rect 680 1158 689 1169
rect 680 1024 689 1076
rect 95 927 104 1020
rect 166 927 175 1015
rect 237 927 246 1015
rect 314 927 323 1016
rect 357 927 366 1016
rect 393 927 402 1013
rect 429 927 438 1013
rect 529 927 538 1013
rect 95 224 104 829
rect 166 722 175 829
rect 166 330 175 624
rect 237 403 246 829
rect 314 722 323 829
rect 166 224 175 276
rect 237 224 246 382
rect 314 370 323 624
rect 314 330 323 349
rect 314 224 323 276
rect 357 224 366 829
rect 393 783 402 829
rect 393 224 402 762
rect 429 757 438 829
rect 529 811 538 829
rect 536 790 538 811
rect 429 224 438 736
rect 529 257 538 790
rect 680 343 689 942
rect 718 709 727 1200
rect 756 1158 765 1169
rect 929 1164 938 1175
rect 756 849 765 1076
rect 842 1024 851 1035
rect 889 1024 898 1111
rect 794 849 803 972
rect 842 849 851 942
rect 889 849 898 942
rect 929 882 938 1082
rect 756 709 765 767
rect 794 709 803 767
rect 842 676 851 767
rect 889 709 898 767
rect 718 556 727 627
rect 756 556 765 627
rect 794 556 803 627
rect 842 540 851 655
rect 889 556 898 627
rect 718 491 727 502
rect 756 453 765 502
rect 794 453 803 502
rect 842 453 851 519
rect 889 453 898 502
rect 929 453 938 861
rect 1005 849 1014 860
rect 967 709 976 828
rect 1005 676 1014 767
rect 967 590 976 627
rect 1005 590 1014 655
rect 1013 569 1014 590
rect 967 556 976 569
rect 1005 540 1014 569
rect 680 253 689 289
rect 529 224 538 236
rect 95 61 104 170
rect 166 147 175 170
rect 166 90 175 126
rect 237 118 246 170
rect 314 118 323 170
rect 357 118 366 170
rect 393 118 402 170
rect 429 154 438 170
rect 529 150 538 170
rect 680 117 689 199
rect 756 88 765 399
rect 794 327 803 399
rect 842 343 851 399
rect 889 343 898 399
rect 794 231 803 306
rect 842 278 851 289
rect 889 214 898 289
rect 929 231 938 432
rect 967 411 976 502
rect 1005 444 1014 519
rect 1005 379 1014 390
rect 794 166 803 177
rect 929 166 938 177
<< ndiffusion >>
rect 163 276 166 330
rect 175 276 178 330
rect 311 276 314 330
rect 323 276 331 330
rect 715 502 718 556
rect 727 502 756 556
rect 765 502 794 556
rect 803 502 806 556
rect 886 502 889 556
rect 898 502 901 556
rect 964 502 967 556
rect 976 502 979 556
rect 753 399 756 453
rect 765 399 794 453
rect 803 399 811 453
rect 832 399 842 453
rect 851 399 889 453
rect 898 399 901 453
rect 677 289 680 343
rect 689 289 692 343
rect 92 170 95 224
rect 104 170 166 224
rect 175 170 212 224
rect 233 170 237 224
rect 246 170 314 224
rect 323 170 333 224
rect 354 170 357 224
rect 366 170 369 224
rect 390 170 393 224
rect 402 170 429 224
rect 438 170 441 224
rect 526 170 529 224
rect 538 170 541 224
rect 677 199 680 253
rect 689 199 692 253
rect 832 289 842 343
rect 851 289 889 343
rect 898 289 901 343
rect 791 177 794 231
rect 803 177 806 231
rect 1002 390 1005 444
rect 1014 390 1017 444
rect 926 177 929 231
rect 938 177 941 231
<< pdiffusion >>
rect 677 1076 680 1158
rect 689 1076 692 1158
rect 677 942 680 1024
rect 689 942 692 1024
rect 92 829 95 927
rect 104 829 113 927
rect 134 829 166 927
rect 175 829 192 927
rect 213 829 237 927
rect 246 829 254 927
rect 275 829 314 927
rect 323 829 333 927
rect 354 829 357 927
rect 366 829 369 927
rect 390 829 393 927
rect 402 829 405 927
rect 426 829 429 927
rect 438 829 441 927
rect 526 829 529 927
rect 538 829 541 927
rect 163 624 166 722
rect 175 624 178 722
rect 311 624 314 722
rect 323 624 331 722
rect 753 1076 756 1158
rect 765 1076 768 1158
rect 926 1082 929 1164
rect 938 1082 941 1164
rect 833 942 842 1024
rect 851 942 859 1024
rect 880 942 889 1024
rect 898 942 903 1024
rect 753 767 756 849
rect 765 767 768 849
rect 789 767 794 849
rect 803 767 812 849
rect 833 767 842 849
rect 851 767 865 849
rect 886 767 889 849
rect 898 767 903 849
rect 715 627 718 709
rect 727 627 732 709
rect 753 627 756 709
rect 765 627 769 709
rect 790 627 794 709
rect 803 627 806 709
rect 886 627 889 709
rect 898 627 903 709
rect 1002 767 1005 849
rect 1014 767 1017 849
rect 964 627 967 709
rect 976 627 979 709
<< ntransistor >>
rect 166 276 175 330
rect 314 276 323 330
rect 718 502 727 556
rect 756 502 765 556
rect 794 502 803 556
rect 889 502 898 556
rect 967 502 976 556
rect 756 399 765 453
rect 794 399 803 453
rect 842 399 851 453
rect 889 399 898 453
rect 680 289 689 343
rect 95 170 104 224
rect 166 170 175 224
rect 237 170 246 224
rect 314 170 323 224
rect 357 170 366 224
rect 393 170 402 224
rect 429 170 438 224
rect 529 170 538 224
rect 680 199 689 253
rect 842 289 851 343
rect 889 289 898 343
rect 794 177 803 231
rect 1005 390 1014 444
rect 929 177 938 231
<< ptransistor >>
rect 680 1076 689 1158
rect 680 942 689 1024
rect 95 829 104 927
rect 166 829 175 927
rect 237 829 246 927
rect 314 829 323 927
rect 357 829 366 927
rect 393 829 402 927
rect 429 829 438 927
rect 529 829 538 927
rect 166 624 175 722
rect 314 624 323 722
rect 756 1076 765 1158
rect 929 1082 938 1164
rect 842 942 851 1024
rect 889 942 898 1024
rect 756 767 765 849
rect 794 767 803 849
rect 842 767 851 849
rect 889 767 898 849
rect 718 627 727 709
rect 756 627 765 709
rect 794 627 803 709
rect 889 627 898 709
rect 1005 767 1014 849
rect 967 627 976 709
<< polycontact >>
rect 712 1200 733 1221
rect 74 749 95 770
rect 225 382 246 403
rect 302 349 323 370
rect 336 352 357 373
rect 381 762 402 783
rect 515 790 536 811
rect 428 736 449 757
rect 879 1111 900 1132
rect 786 972 807 993
rect 918 861 939 882
rect 832 655 853 676
rect 832 519 853 540
rect 955 828 976 849
rect 1005 655 1026 676
rect 956 569 977 590
rect 992 569 1013 590
rect 1005 519 1026 540
rect 927 432 948 453
rect 517 236 538 257
rect 154 126 175 147
rect 674 96 695 117
rect 782 306 803 327
rect 955 390 976 411
rect 879 193 900 214
rect 750 67 771 88
<< ndiffcontact >>
rect 142 276 163 330
rect 178 276 199 330
rect 290 276 311 330
rect 331 276 352 330
rect 694 502 715 556
rect 806 502 827 556
rect 865 502 886 556
rect 901 502 922 556
rect 943 502 964 556
rect 979 502 1000 556
rect 732 399 753 453
rect 811 399 832 453
rect 901 399 922 453
rect 656 289 677 343
rect 692 289 713 343
rect 71 170 92 224
rect 212 170 233 224
rect 333 170 354 224
rect 369 170 390 224
rect 441 170 462 224
rect 505 170 526 224
rect 541 170 562 224
rect 656 199 677 253
rect 692 199 713 253
rect 811 289 832 343
rect 901 289 922 343
rect 770 177 791 231
rect 806 177 827 231
rect 981 390 1002 444
rect 1017 390 1038 444
rect 905 177 926 231
rect 941 177 962 231
<< pdiffcontact >>
rect 656 1076 677 1158
rect 692 1076 713 1158
rect 656 942 677 1024
rect 692 942 713 1024
rect 71 829 92 927
rect 113 829 134 927
rect 192 829 213 927
rect 254 829 275 927
rect 333 829 354 927
rect 369 829 390 927
rect 405 829 426 927
rect 441 829 462 927
rect 505 829 526 927
rect 541 829 562 927
rect 142 624 163 722
rect 178 624 199 722
rect 290 624 311 722
rect 331 624 352 722
rect 732 1076 753 1158
rect 768 1076 789 1158
rect 905 1082 926 1164
rect 941 1082 962 1164
rect 812 942 833 1024
rect 859 942 880 1024
rect 903 942 924 1024
rect 732 767 753 849
rect 768 767 789 849
rect 812 767 833 849
rect 865 767 886 849
rect 903 767 924 849
rect 694 627 715 709
rect 732 627 753 709
rect 769 627 790 709
rect 806 627 827 709
rect 865 627 886 709
rect 903 627 924 709
rect 981 767 1002 849
rect 1017 767 1038 849
rect 943 627 964 709
rect 979 627 1000 709
<< psubstratetap >>
rect 51 30 890 51
<< nsubstratetap >>
rect 42 1292 950 1313
<< metal1 >>
rect 0 1313 1056 1324
rect 0 1292 42 1313
rect 950 1292 1056 1313
rect 0 1284 644 1292
rect 663 1284 1056 1292
rect 0 1260 214 1272
rect 0 1233 67 1245
rect 260 1008 272 1284
rect 324 1260 1056 1272
rect 477 1233 990 1245
rect 260 973 272 989
rect 75 963 207 972
rect 75 960 192 963
rect 75 927 87 960
rect 260 961 304 973
rect 195 927 207 944
rect 260 927 272 961
rect 292 848 304 961
rect 375 952 458 964
rect 339 927 351 944
rect 375 927 387 952
rect 446 927 458 952
rect 477 864 489 1233
rect 1009 1233 1056 1245
rect 541 1205 712 1217
rect 508 927 520 987
rect 541 927 553 1205
rect 701 1170 780 1182
rect 644 1059 656 1170
rect 701 1158 713 1170
rect 768 1158 780 1170
rect 789 1115 879 1127
rect 900 1111 905 1132
rect 732 1059 744 1076
rect 941 1059 953 1082
rect 644 1047 953 1059
rect 121 817 133 829
rect 409 817 421 829
rect 121 805 421 817
rect 446 806 458 829
rect 550 815 562 829
rect 446 794 515 806
rect 549 803 562 815
rect 50 753 74 765
rect 47 349 83 361
rect 47 141 59 349
rect 80 224 92 236
rect 114 145 126 774
rect 147 766 381 778
rect 147 722 159 766
rect 449 740 474 752
rect 296 722 308 734
rect 199 670 290 682
rect 143 330 155 624
rect 213 386 225 398
rect 336 373 348 624
rect 287 354 302 366
rect 336 330 348 352
rect 199 282 290 326
rect 181 248 193 276
rect 181 236 227 248
rect 215 224 227 236
rect 341 240 517 252
rect 215 158 227 170
rect 267 158 279 234
rect 341 224 353 240
rect 550 224 562 803
rect 644 744 656 1047
rect 859 1024 871 1047
rect 713 976 786 988
rect 807 972 812 993
rect 821 930 833 942
rect 907 930 919 942
rect 821 918 919 930
rect 777 894 963 906
rect 777 849 789 894
rect 874 861 918 873
rect 874 849 886 861
rect 951 849 963 894
rect 951 828 955 849
rect 976 828 981 849
rect 732 744 744 767
rect 812 744 824 767
rect 903 744 915 767
rect 1017 744 1029 767
rect 644 732 1029 744
rect 694 709 706 732
rect 769 709 781 732
rect 865 709 877 732
rect 943 709 955 732
rect 827 655 832 676
rect 1000 655 1005 676
rect 741 615 753 627
rect 806 615 818 627
rect 741 603 818 615
rect 912 615 924 627
rect 979 615 991 627
rect 912 603 991 615
rect 955 590 978 591
rect 955 569 956 590
rect 977 569 978 590
rect 955 568 978 569
rect 991 590 1014 591
rect 991 569 992 590
rect 1013 569 1014 590
rect 991 568 1014 569
rect 827 519 832 540
rect 922 522 943 534
rect 1000 519 1005 540
rect 694 490 706 502
rect 865 490 877 502
rect 644 478 877 490
rect 462 187 505 199
rect 369 158 381 170
rect 450 158 462 170
rect 0 129 59 141
rect 128 131 154 143
rect 267 146 381 158
rect 580 141 592 382
rect 644 172 656 478
rect 811 453 823 478
rect 922 432 927 453
rect 741 378 753 399
rect 976 390 981 411
rect 1017 378 1029 390
rect 741 366 1029 378
rect 803 306 811 327
rect 701 277 713 289
rect 901 277 913 289
rect 701 265 913 277
rect 713 219 770 231
rect 900 193 905 214
rect 815 165 827 177
rect 941 165 953 177
rect 815 153 953 165
rect 580 129 1056 141
rect 0 100 674 112
rect 695 100 1056 112
rect 0 71 750 83
rect 771 71 1056 83
rect 0 52 644 55
rect 0 51 450 52
rect 469 51 644 52
rect 663 51 1056 55
rect 0 30 51 51
rect 890 30 1056 51
rect 0 23 210 30
rect 229 23 1056 30
rect 0 15 1056 23
<< m2contact >>
rect 644 1292 663 1303
rect 644 1284 663 1292
rect 214 1253 233 1272
rect 67 1229 86 1248
rect 305 1253 324 1272
rect 257 989 276 1008
rect 192 944 211 963
rect 334 944 353 963
rect 291 829 310 848
rect 990 1229 1009 1248
rect 502 987 521 1006
rect 644 1170 663 1189
rect 474 845 493 864
rect 110 774 129 793
rect 31 753 50 772
rect 83 349 102 368
rect 77 236 96 255
rect 293 734 312 753
rect 474 740 493 759
rect 194 383 213 402
rect 268 351 287 370
rect 263 234 282 253
rect 957 570 976 589
rect 993 570 1012 589
rect 575 382 594 401
rect 109 126 128 145
rect 212 139 231 158
rect 447 139 466 158
rect 644 153 663 172
rect 450 51 469 52
rect 644 51 663 55
rect 210 30 229 42
rect 450 33 469 51
rect 644 36 663 51
rect 210 23 229 30
<< metal2 >>
rect 33 772 47 1339
rect 99 1330 113 1339
rect 99 1316 124 1330
rect 33 0 47 753
rect 68 397 82 1229
rect 110 793 124 1316
rect 233 1257 305 1271
rect 644 1189 658 1284
rect 276 989 502 1003
rect 211 946 334 960
rect 293 753 307 829
rect 476 759 490 845
rect 957 590 971 1339
rect 990 1248 1004 1339
rect 957 589 973 590
rect 990 589 1004 1229
rect 990 570 993 589
rect 957 569 973 570
rect 68 383 194 397
rect 271 384 575 398
rect 271 370 285 384
rect 102 351 268 365
rect 96 237 263 251
rect 110 25 124 126
rect 212 42 226 139
rect 452 52 466 139
rect 644 55 658 153
rect 99 11 124 25
rect 99 0 113 11
rect 957 0 971 569
rect 990 0 1004 570
<< labels >>
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal2 33 0 47 0 1 D
rlabel metal2 99 0 113 0 1 Load
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 SDI
rlabel metal2 99 1339 113 1339 5 Load
rlabel metal2 33 1339 47 1339 5 D
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 1056 1284 1056 1324 7 Vdd!
rlabel metal1 1056 1260 1056 1272 7 ScanReturn
rlabel metal1 1056 129 1056 141 1 Test
rlabel metal1 1056 100 1056 112 1 Clock
rlabel metal1 1056 71 1056 83 1 nReset
rlabel metal1 1056 15 1056 55 1 GND!
rlabel metal1 1056 1233 1056 1245 7 Q
rlabel metal2 957 0 971 0 1 nQ
rlabel metal2 957 1339 971 1339 5 nQ
rlabel metal2 990 0 1004 0 1 Q
rlabel metal2 990 1339 1004 1339 5 Q
<< end >>
