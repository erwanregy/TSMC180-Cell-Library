magic
tech tsmc180
timestamp 1701690570
<< nwell >>
rect 0 605 297 1324
<< polysilicon >>
rect 83 780 92 798
rect 121 780 130 798
rect 158 780 167 798
rect 195 780 204 798
rect 83 620 92 682
rect 121 618 130 682
rect 158 623 167 682
rect 83 566 92 599
rect 195 622 204 682
rect 121 566 130 597
rect 158 566 167 602
rect 195 566 204 601
rect 83 501 92 512
rect 121 501 130 512
rect 158 501 167 512
rect 195 501 204 512
<< ndiffusion >>
rect 80 512 83 566
rect 92 512 121 566
rect 130 512 158 566
rect 167 512 195 566
rect 204 512 207 566
<< pdiffusion >>
rect 80 682 83 780
rect 92 682 96 780
rect 118 682 121 780
rect 130 682 133 780
rect 155 682 158 780
rect 167 682 170 780
rect 192 682 195 780
rect 204 682 207 780
<< nohmic >>
rect 117 1285 152 1286
<< ntransistor >>
rect 83 512 92 566
rect 121 512 130 566
rect 158 512 167 566
rect 195 512 204 566
<< ptransistor >>
rect 83 682 92 780
rect 121 682 130 780
rect 158 682 167 780
rect 195 682 204 780
<< polycontact >>
rect 77 599 98 620
rect 115 597 136 618
rect 152 602 173 623
rect 189 601 210 622
<< ndiffcontact >>
rect 59 512 80 566
rect 207 512 228 566
<< pdiffcontact >>
rect 58 682 80 780
rect 96 682 118 780
rect 133 682 155 780
rect 170 682 192 780
rect 207 682 229 780
<< psubstratetap >>
rect 188 17 223 52
<< nsubstratetap >>
rect 117 1286 152 1320
<< metal1 >>
rect 0 1320 297 1324
rect 0 1314 117 1320
rect 0 1295 39 1314
rect 58 1295 117 1314
rect 0 1286 117 1295
rect 152 1286 297 1320
rect 0 1284 297 1286
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 37 1153 59 1191
rect 37 1131 80 1153
rect 58 868 80 1131
rect 58 846 229 868
rect 58 780 80 846
rect 133 780 155 846
rect 207 780 229 846
rect 102 648 114 682
rect 174 648 186 682
rect 102 636 236 648
rect 151 623 174 624
rect 76 620 99 621
rect 76 599 77 620
rect 98 599 99 620
rect 76 598 99 599
rect 114 618 137 619
rect 114 597 115 618
rect 136 597 137 618
rect 151 602 152 623
rect 173 602 174 623
rect 151 601 174 602
rect 188 622 211 623
rect 188 601 189 622
rect 210 601 211 622
rect 188 600 211 601
rect 224 617 236 636
rect 224 605 259 617
rect 114 596 137 597
rect 224 588 236 605
rect 216 576 236 588
rect 216 566 228 576
rect 59 186 80 512
rect 59 167 60 186
rect 79 167 80 186
rect 59 166 80 167
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 52 297 55
rect 0 47 188 52
rect 0 28 60 47
rect 79 28 188 47
rect 0 17 188 28
rect 223 17 297 52
rect 0 15 297 17
<< m2contact >>
rect 39 1295 58 1314
rect 38 1191 60 1213
rect 77 599 98 620
rect 115 597 136 618
rect 152 602 173 623
rect 189 601 210 622
rect 259 602 278 621
rect 60 167 79 186
rect 60 28 79 47
<< metal2 >>
rect 41 1213 55 1295
rect 99 973 113 1339
rect 81 959 113 973
rect 81 620 95 959
rect 132 945 146 1339
rect 119 931 146 945
rect 119 618 133 931
rect 165 917 179 1339
rect 156 903 179 917
rect 156 623 170 903
rect 198 895 212 1339
rect 193 880 212 895
rect 193 702 207 880
rect 193 688 212 702
rect 80 383 94 599
rect 193 622 207 688
rect 119 411 133 597
rect 156 439 170 602
rect 264 621 278 1339
rect 193 468 207 601
rect 193 454 212 468
rect 156 425 179 439
rect 119 397 146 411
rect 80 369 113 383
rect 62 47 76 167
rect 99 0 113 369
rect 132 0 146 397
rect 165 0 179 425
rect 198 0 212 454
rect 264 0 278 602
<< labels >>
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal2 132 1339 146 1339 5 B
rlabel metal2 165 1339 179 1339 5 C
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal2 165 0 179 0 1 C
rlabel metal2 132 0 146 0 1 B
rlabel metal2 99 0 113 0 1 A
rlabel metal2 198 1339 212 1339 5 D
rlabel metal2 99 1339 113 1339 5 A
rlabel metal2 198 0 212 0 1 D
rlabel metal2 264 0 278 0 1 Y
rlabel metal2 264 1339 278 1339 5 Y
<< end >>
