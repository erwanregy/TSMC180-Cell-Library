magic
tech tsmc180
timestamp 1701546327
<< nwell >>
rect 0 605 627 1328
<< polysilicon >>
rect 95 927 104 1020
rect 166 927 175 1015
rect 237 927 246 1015
rect 314 927 323 1016
rect 357 927 366 1016
rect 393 927 402 1013
rect 429 927 438 1013
rect 529 927 538 1013
rect 95 224 104 829
rect 166 722 175 829
rect 166 330 175 624
rect 237 403 246 829
rect 314 722 323 829
rect 166 224 175 276
rect 237 224 246 382
rect 314 370 323 624
rect 314 330 323 349
rect 314 224 323 276
rect 357 224 366 829
rect 393 783 402 829
rect 393 224 402 762
rect 429 757 438 829
rect 529 811 538 829
rect 536 790 538 811
rect 429 224 438 736
rect 529 257 538 790
rect 529 224 538 236
rect 95 61 104 170
rect 166 147 175 170
rect 166 58 175 126
rect 237 118 246 170
rect 314 118 323 170
rect 357 118 366 170
rect 393 118 402 170
rect 429 154 438 170
rect 529 150 538 170
<< ndiffusion >>
rect 163 276 166 330
rect 175 276 178 330
rect 311 276 314 330
rect 323 276 331 330
rect 92 170 95 224
rect 104 170 166 224
rect 175 170 212 224
rect 233 170 237 224
rect 246 170 314 224
rect 323 170 333 224
rect 354 170 357 224
rect 366 170 369 224
rect 390 170 393 224
rect 402 170 429 224
rect 438 170 441 224
rect 526 170 529 224
rect 538 170 541 224
<< pdiffusion >>
rect 92 829 95 927
rect 104 829 113 927
rect 134 829 166 927
rect 175 829 192 927
rect 213 829 237 927
rect 246 829 254 927
rect 275 829 314 927
rect 323 829 333 927
rect 354 829 357 927
rect 366 829 369 927
rect 390 829 393 927
rect 402 829 405 927
rect 426 829 429 927
rect 438 829 441 927
rect 526 829 529 927
rect 538 829 541 927
rect 163 624 166 722
rect 175 624 178 722
rect 311 624 314 722
rect 323 624 331 722
<< pohmic >>
rect 427 19 430 55
<< ntransistor >>
rect 166 276 175 330
rect 314 276 323 330
rect 95 170 104 224
rect 166 170 175 224
rect 237 170 246 224
rect 314 170 323 224
rect 357 170 366 224
rect 393 170 402 224
rect 429 170 438 224
rect 529 170 538 224
<< ptransistor >>
rect 95 829 104 927
rect 166 829 175 927
rect 237 829 246 927
rect 314 829 323 927
rect 357 829 366 927
rect 393 829 402 927
rect 429 829 438 927
rect 529 829 538 927
rect 166 624 175 722
rect 314 624 323 722
<< polycontact >>
rect 74 749 95 770
rect 225 382 246 403
rect 302 349 323 370
rect 336 352 357 373
rect 381 762 402 783
rect 515 790 536 811
rect 428 736 449 757
rect 517 236 538 257
rect 154 126 175 147
<< ndiffcontact >>
rect 142 276 163 330
rect 178 276 199 330
rect 290 276 311 330
rect 331 276 352 330
rect 71 170 92 224
rect 212 170 233 224
rect 333 170 354 224
rect 369 170 390 224
rect 441 170 462 224
rect 505 170 526 224
rect 541 170 562 224
<< pdiffcontact >>
rect 71 829 92 927
rect 113 829 134 927
rect 192 829 213 927
rect 254 829 275 927
rect 333 829 354 927
rect 369 829 390 927
rect 405 829 426 927
rect 441 829 462 927
rect 505 829 526 927
rect 541 829 562 927
rect 142 624 163 722
rect 178 624 199 722
rect 290 624 311 722
rect 331 624 352 722
<< psubstratetap >>
rect 252 19 427 55
<< nsubstratetap >>
rect 136 1293 503 1321
<< metal1 >>
rect 0 1321 627 1328
rect 0 1293 136 1321
rect 503 1293 627 1321
rect 0 1284 627 1293
rect 0 1260 214 1272
rect 0 1233 67 1245
rect 260 1008 272 1284
rect 324 1260 627 1272
rect 477 1233 627 1245
rect 260 973 272 989
rect 75 963 207 972
rect 75 960 192 963
rect 75 927 87 960
rect 260 961 304 973
rect 195 927 207 944
rect 260 927 272 961
rect 292 848 304 961
rect 375 952 458 964
rect 339 927 351 944
rect 375 927 387 952
rect 446 927 458 952
rect 477 864 489 1233
rect 541 1205 627 1217
rect 508 927 520 987
rect 541 927 553 1205
rect 121 817 133 829
rect 409 817 421 829
rect 121 805 421 817
rect 446 806 458 829
rect 550 815 562 829
rect 446 794 515 806
rect 549 803 562 815
rect 50 753 74 765
rect 47 349 83 361
rect 47 141 59 349
rect 80 224 92 236
rect 114 145 126 774
rect 147 766 381 778
rect 147 722 159 766
rect 449 740 474 752
rect 296 722 308 734
rect 199 670 290 682
rect 143 330 155 624
rect 213 386 225 398
rect 336 373 348 624
rect 287 354 302 366
rect 336 330 348 352
rect 199 282 290 326
rect 181 248 193 276
rect 181 236 227 248
rect 215 224 227 236
rect 341 240 517 252
rect 215 158 227 170
rect 267 158 279 234
rect 341 224 353 240
rect 550 224 562 803
rect 462 187 505 199
rect 369 158 381 170
rect 450 158 462 170
rect 0 129 59 141
rect 128 131 154 143
rect 267 146 381 158
rect 580 141 592 382
rect 580 129 627 141
rect 0 100 627 112
rect 0 71 627 83
rect 0 55 627 59
rect 0 42 252 55
rect 0 23 210 42
rect 229 23 252 42
rect 0 19 252 23
rect 427 52 627 55
rect 427 33 450 52
rect 469 33 627 52
rect 427 19 627 33
rect 0 15 627 19
<< m2contact >>
rect 214 1253 233 1272
rect 67 1229 86 1248
rect 305 1253 324 1272
rect 257 989 276 1008
rect 192 944 211 963
rect 334 944 353 963
rect 291 829 310 848
rect 502 987 521 1006
rect 474 845 493 864
rect 110 774 129 793
rect 31 753 50 772
rect 83 349 102 368
rect 77 236 96 255
rect 293 734 312 753
rect 474 740 493 759
rect 194 383 213 402
rect 268 351 287 370
rect 263 234 282 253
rect 575 382 594 401
rect 109 126 128 145
rect 212 139 231 158
rect 447 139 466 158
rect 210 23 229 42
rect 450 33 469 52
<< metal2 >>
rect 33 772 47 1339
rect 99 1330 113 1339
rect 99 1316 124 1330
rect 33 0 47 753
rect 68 397 82 1229
rect 110 793 124 1316
rect 233 1257 305 1271
rect 276 989 502 1003
rect 211 946 334 960
rect 293 753 307 829
rect 476 759 490 845
rect 68 383 194 397
rect 271 384 575 398
rect 271 370 285 384
rect 102 351 268 365
rect 96 237 263 251
rect 110 25 124 126
rect 212 42 226 139
rect 452 52 466 139
rect 99 11 124 25
rect 99 0 113 11
<< labels >>
rlabel metal1 0 1284 0 1328 3 Vdd!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal2 33 0 47 0 1 D
rlabel metal2 99 0 113 0 1 Load
rlabel metal1 0 15 0 59 3 GND!
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 SDI
rlabel metal1 627 1205 627 1217 7 M
rlabel metal1 627 1233 627 1245 7 Q
rlabel metal1 627 1284 627 1328 7 Vdd!
rlabel metal1 627 1260 627 1272 7 ScanReturn
rlabel metal1 627 129 627 141 7 Test
rlabel metal1 627 100 627 112 7 Clock
rlabel metal1 627 71 627 83 7 nReset
rlabel metal1 627 15 627 59 7 GND!
rlabel metal2 99 1339 113 1339 5 Load
rlabel metal2 33 1339 47 1339 5 D
<< end >>
