magic
tech tsmc180
timestamp 1701442775
<< nwell >>
rect 0 632 297 1284
<< polysilicon >>
rect 119 733 128 744
rect 119 623 128 634
rect 119 590 128 602
rect 119 525 128 536
<< ndiffusion >>
rect 116 569 119 590
rect 95 536 119 569
rect 128 557 152 590
rect 128 536 131 557
<< pdiffusion >>
rect 115 712 119 733
rect 94 634 119 712
rect 128 712 134 733
rect 128 634 155 712
<< ntransistor >>
rect 119 536 128 590
<< ptransistor >>
rect 119 634 128 733
<< polycontact >>
rect 108 602 129 623
<< ndiffcontact >>
rect 95 569 116 590
rect 131 536 152 557
<< pdiffcontact >>
rect 94 712 115 733
rect 134 712 155 733
<< psubstratetap >>
rect 169 17 204 52
<< nsubstratetap >>
rect 186 1287 221 1322
<< metal1 >>
rect 0 1322 297 1324
rect 0 1305 186 1322
rect 0 1284 94 1305
rect 115 1287 186 1305
rect 221 1287 297 1322
rect 115 1284 297 1287
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 95 602 108 623
rect 95 590 116 602
rect 152 536 241 557
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 52 241 55
rect 0 17 169 52
rect 204 35 241 52
rect 262 35 297 55
rect 204 17 297 35
rect 0 15 297 17
<< m2contact >>
rect 94 1284 115 1305
rect 94 712 115 733
rect 241 536 262 557
rect 241 35 262 55
<< metal2 >>
rect 132 1305 146 1339
rect 132 1284 155 1305
rect 94 733 115 1284
rect 135 55 155 1284
rect 132 34 155 55
rect 241 55 262 536
rect 132 0 146 34
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal2 132 0 146 0 1 High
rlabel metal2 132 1339 146 1339 5 High
<< end >>