magic
tech tsmc180
timestamp 1701621919
<< nwell >>
rect 545 605 2574 1324
<< polysilicon >>
rect 1107 1172 1116 1183
rect 1147 1172 1156 1183
rect 1187 1172 1196 1183
rect 1227 1172 1236 1183
rect 912 824 921 835
rect 952 824 961 835
rect 992 824 1001 835
rect 1032 824 1041 835
rect 798 772 807 784
rect 836 772 845 784
rect 725 733 734 747
rect 613 719 622 733
rect 613 564 622 621
rect 613 342 622 543
rect 725 529 734 621
rect 798 527 807 621
rect 725 342 734 508
rect 798 361 807 506
rect 836 361 845 621
rect 1709 1170 1718 1181
rect 1749 1170 1758 1181
rect 1789 1170 1798 1181
rect 1829 1170 1838 1181
rect 1514 824 1523 835
rect 1554 824 1563 835
rect 1594 824 1603 835
rect 1634 824 1643 835
rect 1400 772 1409 784
rect 1438 772 1447 784
rect 1327 733 1336 747
rect 912 525 921 620
rect 798 352 845 361
rect 798 342 807 352
rect 836 342 845 352
rect 912 365 921 504
rect 952 365 961 620
rect 992 365 1001 620
rect 1032 365 1041 620
rect 1107 524 1116 621
rect 912 356 1041 365
rect 912 342 921 356
rect 952 342 961 356
rect 992 342 1001 356
rect 1032 342 1041 356
rect 1107 366 1116 503
rect 1147 366 1156 621
rect 1187 366 1196 621
rect 1227 366 1236 621
rect 1327 477 1336 621
rect 1400 477 1409 621
rect 1107 357 1236 366
rect 1107 342 1116 357
rect 1147 342 1156 357
rect 1187 342 1196 357
rect 1227 342 1236 357
rect 1327 342 1336 456
rect 1400 361 1409 456
rect 1438 361 1447 621
rect 1514 477 1523 620
rect 1400 352 1447 361
rect 1400 342 1409 352
rect 1438 342 1447 352
rect 1514 364 1523 456
rect 1554 364 1563 620
rect 1594 364 1603 620
rect 1634 364 1643 620
rect 2315 1168 2324 1179
rect 2355 1168 2364 1179
rect 2395 1168 2404 1179
rect 2435 1168 2444 1179
rect 2120 822 2129 833
rect 2160 822 2169 833
rect 2200 822 2209 833
rect 2240 822 2249 833
rect 2006 770 2015 782
rect 2044 770 2053 782
rect 1933 731 1942 745
rect 1709 478 1718 619
rect 1514 355 1643 364
rect 1514 342 1523 355
rect 1554 342 1563 355
rect 1594 342 1603 355
rect 1634 342 1643 355
rect 1709 371 1718 457
rect 1749 371 1758 619
rect 1789 371 1798 619
rect 1829 371 1838 619
rect 1933 436 1942 619
rect 2006 436 2015 619
rect 1709 362 1838 371
rect 1709 342 1718 362
rect 1749 342 1758 362
rect 1789 342 1798 362
rect 1829 342 1838 362
rect 1933 342 1942 415
rect 2006 361 2015 415
rect 2044 361 2053 619
rect 2120 434 2129 618
rect 2006 352 2053 361
rect 2006 342 2015 352
rect 2044 342 2053 352
rect 2120 364 2129 413
rect 2160 364 2169 618
rect 2200 364 2209 618
rect 2240 364 2249 618
rect 2315 433 2324 617
rect 2120 355 2249 364
rect 2120 342 2129 355
rect 2160 342 2169 355
rect 2200 342 2209 355
rect 2240 342 2249 355
rect 2315 365 2324 412
rect 2355 365 2364 617
rect 2395 365 2404 617
rect 2435 365 2444 617
rect 2315 356 2444 365
rect 2315 342 2324 356
rect 2355 342 2364 356
rect 2395 342 2404 356
rect 2435 342 2444 356
rect 725 289 734 300
rect 613 277 622 288
rect 798 275 807 286
rect 836 275 845 286
rect 912 255 921 266
rect 952 255 961 266
rect 992 255 1001 266
rect 1032 255 1041 266
rect 1327 289 1336 300
rect 1400 275 1409 286
rect 1438 275 1447 286
rect 1514 255 1523 266
rect 1554 255 1563 266
rect 1594 255 1603 266
rect 1634 255 1643 266
rect 1933 289 1942 300
rect 2006 275 2015 286
rect 2044 275 2053 286
rect 2120 255 2129 266
rect 2160 255 2169 266
rect 2200 255 2209 266
rect 2240 255 2249 266
rect 1107 123 1116 135
rect 1147 123 1156 135
rect 1187 123 1196 135
rect 1227 123 1236 135
rect 1709 123 1718 135
rect 1749 123 1758 135
rect 1789 123 1798 135
rect 1829 123 1838 135
rect 2315 123 2324 135
rect 2355 123 2364 135
rect 2395 123 2404 135
rect 2435 123 2444 135
<< ndiffusion >>
rect 608 288 613 342
rect 622 288 627 342
rect 720 300 725 342
rect 734 300 739 342
rect 795 286 798 342
rect 807 286 811 342
rect 832 286 836 342
rect 845 286 850 342
rect 907 266 912 342
rect 921 266 926 342
rect 947 266 952 342
rect 961 266 966 342
rect 987 266 992 342
rect 1001 266 1006 342
rect 1027 266 1032 342
rect 1041 266 1046 342
rect 1102 135 1107 342
rect 1116 135 1121 342
rect 1142 135 1147 342
rect 1156 135 1161 342
rect 1182 135 1187 342
rect 1196 135 1201 342
rect 1222 135 1227 342
rect 1236 135 1241 342
rect 1322 300 1327 342
rect 1336 300 1341 342
rect 1397 286 1400 342
rect 1409 286 1413 342
rect 1434 286 1438 342
rect 1447 286 1452 342
rect 1509 266 1514 342
rect 1523 266 1528 342
rect 1549 266 1554 342
rect 1563 266 1568 342
rect 1589 266 1594 342
rect 1603 266 1608 342
rect 1629 266 1634 342
rect 1643 266 1648 342
rect 1704 135 1709 342
rect 1718 135 1723 342
rect 1744 135 1749 342
rect 1758 135 1763 342
rect 1784 135 1789 342
rect 1798 135 1803 342
rect 1824 135 1829 342
rect 1838 135 1843 342
rect 1928 300 1933 342
rect 1942 300 1947 342
rect 2003 286 2006 342
rect 2015 286 2019 342
rect 2040 286 2044 342
rect 2053 286 2058 342
rect 2115 266 2120 342
rect 2129 266 2134 342
rect 2155 266 2160 342
rect 2169 266 2174 342
rect 2195 266 2200 342
rect 2209 266 2214 342
rect 2235 266 2240 342
rect 2249 266 2254 342
rect 2310 135 2315 342
rect 2324 135 2329 342
rect 2350 135 2355 342
rect 2364 135 2369 342
rect 2390 135 2395 342
rect 2404 135 2409 342
rect 2430 135 2435 342
rect 2444 135 2449 342
<< pdiffusion >>
rect 608 621 613 719
rect 622 621 627 719
rect 720 621 725 733
rect 734 621 739 733
rect 795 621 798 772
rect 807 621 811 772
rect 832 621 836 772
rect 845 621 851 772
rect 907 620 912 824
rect 921 620 926 824
rect 947 620 952 824
rect 961 620 966 824
rect 987 620 992 824
rect 1001 620 1006 824
rect 1027 620 1032 824
rect 1041 620 1046 824
rect 1102 621 1107 1172
rect 1116 621 1121 1172
rect 1142 621 1147 1172
rect 1156 621 1161 1172
rect 1182 621 1187 1172
rect 1196 621 1201 1172
rect 1222 621 1227 1172
rect 1236 621 1241 1172
rect 1322 621 1327 733
rect 1336 621 1341 733
rect 1397 621 1400 772
rect 1409 621 1413 772
rect 1434 621 1438 772
rect 1447 621 1453 772
rect 1509 620 1514 824
rect 1523 620 1528 824
rect 1549 620 1554 824
rect 1563 620 1568 824
rect 1589 620 1594 824
rect 1603 620 1608 824
rect 1629 620 1634 824
rect 1643 620 1648 824
rect 1704 619 1709 1170
rect 1718 619 1723 1170
rect 1744 619 1749 1170
rect 1758 619 1763 1170
rect 1784 619 1789 1170
rect 1798 619 1803 1170
rect 1824 619 1829 1170
rect 1838 619 1843 1170
rect 1928 619 1933 731
rect 1942 619 1947 731
rect 2003 619 2006 770
rect 2015 619 2019 770
rect 2040 619 2044 770
rect 2053 619 2059 770
rect 2115 618 2120 822
rect 2129 618 2134 822
rect 2155 618 2160 822
rect 2169 618 2174 822
rect 2195 618 2200 822
rect 2209 618 2214 822
rect 2235 618 2240 822
rect 2249 618 2254 822
rect 2310 617 2315 1168
rect 2324 617 2329 1168
rect 2350 617 2355 1168
rect 2364 617 2369 1168
rect 2390 617 2395 1168
rect 2404 617 2409 1168
rect 2430 617 2435 1168
rect 2444 617 2449 1168
<< ntransistor >>
rect 613 288 622 342
rect 725 300 734 342
rect 798 286 807 342
rect 836 286 845 342
rect 912 266 921 342
rect 952 266 961 342
rect 992 266 1001 342
rect 1032 266 1041 342
rect 1107 135 1116 342
rect 1147 135 1156 342
rect 1187 135 1196 342
rect 1227 135 1236 342
rect 1327 300 1336 342
rect 1400 286 1409 342
rect 1438 286 1447 342
rect 1514 266 1523 342
rect 1554 266 1563 342
rect 1594 266 1603 342
rect 1634 266 1643 342
rect 1709 135 1718 342
rect 1749 135 1758 342
rect 1789 135 1798 342
rect 1829 135 1838 342
rect 1933 300 1942 342
rect 2006 286 2015 342
rect 2044 286 2053 342
rect 2120 266 2129 342
rect 2160 266 2169 342
rect 2200 266 2209 342
rect 2240 266 2249 342
rect 2315 135 2324 342
rect 2355 135 2364 342
rect 2395 135 2404 342
rect 2435 135 2444 342
<< ptransistor >>
rect 613 621 622 719
rect 725 621 734 733
rect 798 621 807 772
rect 836 621 845 772
rect 912 620 921 824
rect 952 620 961 824
rect 992 620 1001 824
rect 1032 620 1041 824
rect 1107 621 1116 1172
rect 1147 621 1156 1172
rect 1187 621 1196 1172
rect 1227 621 1236 1172
rect 1327 621 1336 733
rect 1400 621 1409 772
rect 1438 621 1447 772
rect 1514 620 1523 824
rect 1554 620 1563 824
rect 1594 620 1603 824
rect 1634 620 1643 824
rect 1709 619 1718 1170
rect 1749 619 1758 1170
rect 1789 619 1798 1170
rect 1829 619 1838 1170
rect 1933 619 1942 731
rect 2006 619 2015 770
rect 2044 619 2053 770
rect 2120 618 2129 822
rect 2160 618 2169 822
rect 2200 618 2209 822
rect 2240 618 2249 822
rect 2315 617 2324 1168
rect 2355 617 2364 1168
rect 2395 617 2404 1168
rect 2435 617 2444 1168
<< polycontact >>
rect 613 543 634 564
rect 713 508 734 529
rect 785 506 807 527
rect 900 504 921 525
rect 1095 503 1116 524
rect 1315 456 1336 477
rect 1387 456 1409 477
rect 1502 456 1523 477
rect 1697 457 1718 478
rect 1921 415 1942 436
rect 1993 415 2015 436
rect 2108 413 2129 434
rect 2303 412 2324 433
<< ndiffcontact >>
rect 587 288 608 342
rect 627 288 648 342
rect 699 300 720 342
rect 739 300 760 342
rect 774 286 795 342
rect 811 286 832 342
rect 850 286 871 342
rect 886 266 907 342
rect 926 266 947 342
rect 966 266 987 342
rect 1006 266 1027 342
rect 1046 266 1067 342
rect 1081 135 1102 342
rect 1121 135 1142 342
rect 1161 135 1182 342
rect 1201 135 1222 342
rect 1241 135 1262 342
rect 1301 300 1322 342
rect 1341 300 1362 342
rect 1376 286 1397 342
rect 1413 286 1434 342
rect 1452 286 1473 342
rect 1488 266 1509 342
rect 1528 266 1549 342
rect 1568 266 1589 342
rect 1608 266 1629 342
rect 1648 266 1669 342
rect 1683 135 1704 342
rect 1723 135 1744 342
rect 1763 135 1784 342
rect 1803 135 1824 342
rect 1843 135 1864 342
rect 1907 300 1928 342
rect 1947 300 1968 342
rect 1982 286 2003 342
rect 2019 286 2040 342
rect 2058 286 2079 342
rect 2094 266 2115 342
rect 2134 266 2155 342
rect 2174 266 2195 342
rect 2214 266 2235 342
rect 2254 266 2275 342
rect 2289 135 2310 342
rect 2329 135 2350 342
rect 2369 135 2390 342
rect 2409 135 2430 342
rect 2449 135 2470 342
<< pdiffcontact >>
rect 587 621 608 719
rect 627 621 648 719
rect 699 621 720 733
rect 739 621 760 733
rect 774 621 795 772
rect 811 621 832 772
rect 851 621 872 772
rect 886 620 907 824
rect 926 620 947 824
rect 966 620 987 824
rect 1006 620 1027 824
rect 1046 620 1067 824
rect 1081 621 1102 1172
rect 1121 621 1142 1172
rect 1161 621 1182 1172
rect 1201 621 1222 1172
rect 1241 621 1262 1172
rect 1301 621 1322 733
rect 1341 621 1362 733
rect 1376 621 1397 772
rect 1413 621 1434 772
rect 1453 621 1474 772
rect 1488 620 1509 824
rect 1528 620 1549 824
rect 1568 620 1589 824
rect 1608 620 1629 824
rect 1648 620 1669 824
rect 1683 619 1704 1170
rect 1723 619 1744 1170
rect 1763 619 1784 1170
rect 1803 619 1824 1170
rect 1843 619 1864 1170
rect 1907 619 1928 731
rect 1947 619 1968 731
rect 1982 619 2003 770
rect 2019 619 2040 770
rect 2059 619 2080 770
rect 2094 618 2115 822
rect 2134 618 2155 822
rect 2174 618 2195 822
rect 2214 618 2235 822
rect 2254 618 2275 822
rect 2289 617 2310 1168
rect 2329 617 2350 1168
rect 2369 617 2390 1168
rect 2409 617 2430 1168
rect 2449 617 2470 1168
<< psubstratetap >>
rect 819 18 854 53
rect 876 19 911 54
rect 987 16 1022 51
rect 1177 15 1212 50
rect 1323 15 1358 50
rect 1393 15 1428 50
rect 1606 16 1641 51
rect 1715 15 1750 50
rect 1825 15 1860 50
rect 2071 15 2106 50
rect 2234 16 2269 51
rect 2362 15 2397 50
rect 2436 15 2471 50
rect 2492 15 2527 50
<< nsubstratetap >>
rect 657 1284 692 1319
rect 810 1289 845 1324
rect 1120 1287 1155 1322
rect 1329 1286 1364 1321
rect 1516 1288 1551 1323
rect 1707 1284 1742 1319
rect 1801 1289 1836 1324
rect 2007 1286 2042 1321
rect 2127 1287 2162 1322
rect 2205 1289 2240 1324
rect 2399 1288 2434 1323
rect 2489 1286 2524 1321
<< metal1 >>
rect 219 1319 810 1324
rect 219 1313 657 1319
rect 219 1292 627 1313
rect 648 1292 657 1313
rect 219 1284 657 1292
rect 692 1314 810 1319
rect 692 1313 774 1314
rect 692 1292 699 1313
rect 720 1293 774 1313
rect 795 1293 810 1314
rect 720 1292 810 1293
rect 692 1289 810 1292
rect 845 1323 1801 1324
rect 845 1322 1516 1323
rect 845 1317 1120 1322
rect 845 1296 851 1317
rect 872 1313 1120 1317
rect 872 1312 966 1313
rect 872 1296 886 1312
rect 845 1291 886 1296
rect 907 1292 966 1312
rect 987 1292 1046 1313
rect 1067 1292 1081 1313
rect 1102 1292 1120 1313
rect 907 1291 1120 1292
rect 845 1289 1120 1291
rect 692 1287 1120 1289
rect 1155 1321 1516 1322
rect 1155 1315 1329 1321
rect 1155 1313 1301 1315
rect 1155 1292 1161 1313
rect 1182 1292 1241 1313
rect 1262 1296 1301 1313
rect 1322 1296 1329 1315
rect 1262 1292 1329 1296
rect 1155 1287 1329 1292
rect 692 1286 1329 1287
rect 1364 1313 1516 1321
rect 1364 1309 1488 1313
rect 1364 1290 1376 1309
rect 1397 1290 1453 1309
rect 1474 1294 1488 1309
rect 1509 1294 1516 1313
rect 1474 1290 1516 1294
rect 1364 1288 1516 1290
rect 1551 1319 1801 1323
rect 1551 1314 1707 1319
rect 1551 1313 1683 1314
rect 1551 1310 1648 1313
rect 1551 1291 1568 1310
rect 1589 1294 1648 1310
rect 1669 1295 1683 1313
rect 1704 1295 1707 1314
rect 1669 1294 1707 1295
rect 1589 1291 1707 1294
rect 1551 1288 1707 1291
rect 1364 1286 1707 1288
rect 692 1284 1707 1286
rect 1742 1313 1801 1319
rect 1742 1294 1763 1313
rect 1784 1294 1801 1313
rect 1742 1289 1801 1294
rect 1836 1322 2205 1324
rect 1836 1321 2127 1322
rect 1836 1314 2007 1321
rect 1836 1295 1843 1314
rect 1864 1295 1907 1314
rect 1928 1313 2007 1314
rect 1928 1295 1982 1313
rect 1836 1294 1982 1295
rect 2003 1294 2007 1313
rect 1836 1289 2007 1294
rect 1742 1286 2007 1289
rect 2042 1314 2127 1321
rect 2042 1312 2094 1314
rect 2042 1293 2059 1312
rect 2080 1295 2094 1312
rect 2115 1295 2127 1314
rect 2080 1293 2127 1295
rect 2042 1287 2127 1293
rect 2162 1308 2205 1322
rect 2162 1289 2174 1308
rect 2195 1289 2205 1308
rect 2240 1323 2574 1324
rect 2240 1314 2399 1323
rect 2240 1295 2254 1314
rect 2275 1295 2289 1314
rect 2310 1311 2399 1314
rect 2310 1295 2369 1311
rect 2240 1292 2369 1295
rect 2390 1292 2399 1311
rect 2240 1289 2399 1292
rect 2162 1288 2399 1289
rect 2434 1321 2574 1323
rect 2434 1316 2489 1321
rect 2434 1297 2449 1316
rect 2470 1297 2489 1316
rect 2434 1288 2489 1297
rect 2162 1287 2489 1288
rect 2042 1286 2489 1287
rect 2524 1286 2574 1321
rect 1742 1284 2574 1286
rect 446 1257 557 1269
rect 682 1260 2574 1272
rect 2500 1237 2574 1245
rect 447 1233 2574 1237
rect 447 1225 2512 1233
rect 1081 1172 1102 1189
rect 1161 1172 1182 1189
rect 1241 1172 1262 1189
rect 627 719 648 772
rect 699 733 720 916
rect 774 772 795 916
rect 851 772 872 915
rect 886 824 907 915
rect 966 824 987 915
rect 1046 824 1067 915
rect 587 561 601 621
rect 575 546 601 561
rect 479 515 556 527
rect 512 463 556 475
rect 587 342 601 546
rect 634 547 659 559
rect 659 514 713 526
rect 746 524 760 621
rect 746 509 785 524
rect 746 342 760 509
rect 820 520 832 621
rect 1683 1170 1704 1190
rect 1763 1170 1784 1190
rect 1843 1170 1864 1190
rect 1301 733 1322 916
rect 1376 772 1397 916
rect 1453 772 1474 915
rect 1488 824 1509 915
rect 1568 824 1589 915
rect 1648 824 1669 915
rect 931 608 944 620
rect 1011 608 1023 620
rect 931 595 1023 608
rect 1126 609 1139 621
rect 1206 609 1218 621
rect 1126 596 1257 609
rect 820 508 900 520
rect 820 342 832 508
rect 1010 519 1023 595
rect 1242 524 1257 596
rect 1010 507 1095 519
rect 1010 367 1023 507
rect 1242 509 1269 524
rect 1242 367 1257 509
rect 1288 460 1315 472
rect 1348 474 1362 621
rect 1348 459 1387 474
rect 933 354 1023 367
rect 933 342 946 354
rect 1010 342 1023 354
rect 1128 354 1257 367
rect 1128 342 1141 354
rect 1205 342 1218 354
rect 1348 342 1362 459
rect 1422 472 1434 621
rect 1533 608 1546 620
rect 1613 608 1625 620
rect 2289 1168 2310 1188
rect 2369 1168 2390 1188
rect 2449 1168 2470 1188
rect 1907 731 1928 914
rect 1982 770 2003 914
rect 2059 770 2080 913
rect 2094 822 2115 913
rect 2174 822 2195 913
rect 2254 822 2275 913
rect 1533 595 1625 608
rect 1422 460 1502 472
rect 1422 342 1434 460
rect 1612 473 1625 595
rect 1728 607 1741 619
rect 1808 607 1820 619
rect 1728 594 1859 607
rect 1612 461 1697 473
rect 1612 367 1625 461
rect 1844 477 1859 594
rect 1844 462 1877 477
rect 1844 367 1859 462
rect 1895 419 1921 431
rect 1954 433 1968 619
rect 1954 418 1993 433
rect 1535 354 1625 367
rect 1535 342 1548 354
rect 1612 342 1625 354
rect 1730 354 1859 367
rect 1730 342 1743 354
rect 1807 342 1820 354
rect 1954 342 1968 418
rect 2028 429 2040 619
rect 2139 606 2152 618
rect 2219 606 2231 618
rect 2139 593 2231 606
rect 2028 417 2108 429
rect 2028 342 2040 417
rect 2218 428 2231 593
rect 2334 605 2347 617
rect 2414 605 2426 617
rect 2334 592 2465 605
rect 2218 416 2303 428
rect 2218 367 2231 416
rect 2450 423 2465 592
rect 2450 411 2494 423
rect 2450 367 2465 411
rect 2141 354 2231 367
rect 2141 342 2154 354
rect 2218 342 2231 354
rect 2336 354 2465 367
rect 2336 342 2349 354
rect 2413 342 2426 354
rect 627 277 648 288
rect 626 55 647 277
rect 699 55 720 300
rect 774 55 795 286
rect 850 55 871 286
rect 886 55 907 266
rect 966 55 987 266
rect 1047 55 1064 266
rect 1083 55 1098 135
rect 1164 55 1179 135
rect 1242 134 1258 135
rect 1243 55 1258 134
rect 1301 55 1322 300
rect 1376 55 1397 286
rect 1452 55 1473 286
rect 1490 55 1507 266
rect 1568 55 1589 266
rect 1649 55 1666 266
rect 1685 55 1700 135
rect 1766 55 1781 135
rect 1844 134 1860 135
rect 1845 55 1860 134
rect 1907 55 1928 300
rect 1982 55 2003 286
rect 2058 55 2079 286
rect 2096 55 2113 266
rect 2174 55 2195 266
rect 2255 55 2272 266
rect 2291 55 2306 135
rect 2372 55 2387 135
rect 2450 134 2466 135
rect 2451 55 2466 134
rect 2482 83 2494 411
rect 2506 112 2518 458
rect 2531 141 2543 506
rect 2531 129 2574 141
rect 2506 100 2574 112
rect 2482 71 2574 83
rect 626 54 2574 55
rect 626 53 876 54
rect 626 18 819 53
rect 854 19 876 53
rect 911 51 2574 54
rect 911 19 987 51
rect 854 18 987 19
rect 626 16 987 18
rect 1022 50 1606 51
rect 1022 16 1177 50
rect 626 15 1177 16
rect 1212 15 1323 50
rect 1358 15 1393 50
rect 1428 16 1606 50
rect 1641 50 2234 51
rect 1641 16 1715 50
rect 1428 15 1715 16
rect 1750 15 1825 50
rect 1860 15 2071 50
rect 2106 16 2234 50
rect 2269 50 2574 51
rect 2269 16 2362 50
rect 2106 15 2362 16
rect 2397 15 2436 50
rect 2471 15 2492 50
rect 2527 15 2574 50
<< m2contact >>
rect 179 1284 219 1324
rect 627 1292 648 1313
rect 699 1292 720 1313
rect 774 1293 795 1314
rect 851 1296 872 1317
rect 886 1291 907 1312
rect 966 1292 987 1313
rect 1046 1292 1067 1313
rect 1081 1292 1102 1313
rect 1161 1292 1182 1313
rect 1241 1292 1262 1313
rect 1301 1296 1322 1315
rect 1376 1290 1397 1309
rect 1453 1290 1474 1309
rect 1488 1294 1509 1313
rect 1568 1291 1589 1310
rect 1648 1294 1669 1313
rect 1683 1295 1704 1314
rect 1763 1294 1784 1313
rect 1843 1295 1864 1314
rect 1907 1295 1928 1314
rect 1982 1294 2003 1313
rect 2059 1293 2080 1312
rect 2094 1295 2115 1314
rect 2174 1289 2195 1308
rect 2254 1295 2275 1314
rect 2289 1295 2310 1314
rect 2369 1292 2390 1311
rect 2449 1297 2470 1316
rect 427 1253 446 1272
rect 557 1253 576 1272
rect 663 1253 682 1272
rect 428 1218 447 1237
rect 1081 1189 1102 1210
rect 1161 1189 1182 1210
rect 1241 1189 1262 1210
rect 699 916 720 937
rect 627 772 648 793
rect 774 916 795 937
rect 851 915 872 936
rect 886 915 907 936
rect 966 915 987 936
rect 1046 915 1067 936
rect 556 544 575 563
rect 460 511 479 530
rect 556 511 575 530
rect 493 461 512 480
rect 556 460 575 479
rect 659 544 678 563
rect 640 510 659 529
rect 1683 1190 1704 1211
rect 1763 1190 1784 1211
rect 1843 1190 1864 1211
rect 1301 916 1322 937
rect 1376 916 1397 937
rect 1453 915 1474 936
rect 1488 915 1509 936
rect 1568 915 1589 936
rect 1648 915 1669 936
rect 1269 507 1288 526
rect 1269 457 1288 476
rect 2289 1188 2310 1209
rect 2369 1188 2390 1209
rect 2449 1188 2470 1209
rect 1907 914 1928 935
rect 1982 914 2003 935
rect 2059 913 2080 934
rect 2094 913 2115 934
rect 2174 913 2195 934
rect 2254 913 2275 934
rect 1877 460 1896 479
rect 1876 416 1895 435
rect 2524 506 2543 525
rect 2499 458 2518 477
<< metal2 >>
rect 0 1324 400 1339
rect 0 1284 179 1324
rect 219 1284 400 1324
rect 0 0 400 1284
rect 429 1272 443 1339
rect 429 0 443 1218
rect 462 530 476 1339
rect 462 0 476 511
rect 495 480 509 1339
rect 495 0 509 461
rect 528 432 542 1339
rect 559 563 573 1253
rect 627 793 648 1292
rect 663 563 677 1253
rect 699 937 720 1292
rect 774 937 795 1293
rect 851 936 872 1296
rect 886 936 907 1291
rect 966 936 987 1292
rect 1046 936 1067 1292
rect 1081 1210 1102 1292
rect 1161 1210 1182 1292
rect 1241 1210 1262 1292
rect 1301 937 1322 1296
rect 1376 937 1397 1290
rect 1453 936 1474 1290
rect 1488 936 1509 1294
rect 1568 936 1589 1291
rect 1648 936 1669 1294
rect 1683 1211 1704 1295
rect 1763 1211 1784 1294
rect 1843 1211 1864 1295
rect 1907 935 1928 1295
rect 1982 935 2003 1294
rect 2059 934 2080 1293
rect 2094 934 2115 1295
rect 2174 934 2195 1289
rect 2254 934 2275 1295
rect 2289 1209 2310 1295
rect 2369 1209 2390 1292
rect 2449 1209 2470 1297
rect 575 512 640 526
rect 1288 508 2524 522
rect 575 460 1269 474
rect 1896 460 2499 474
rect 528 418 1876 432
rect 528 0 542 418
<< labels >>
rlabel metal2 0 0 400 0 1 Vdd!
rlabel metal2 462 0 476 0 1 Test
rlabel metal2 495 0 509 0 1 Clock
rlabel metal2 528 0 542 0 1 nReset
rlabel metal2 429 0 443 0 1 SDI
rlabel metal2 0 1339 400 1339 5 Vdd!
rlabel metal2 429 1339 443 1339 5 SDO
rlabel metal2 495 1339 509 1339 5 Clock
rlabel metal2 462 1339 476 1339 5 Test
rlabel metal2 528 1339 542 1339 5 nReset
rlabel metal1 2574 15 2574 55 7 GND!
rlabel metal1 2574 129 2574 141 7 TestOut
rlabel metal1 2574 100 2574 112 7 ClockOut
rlabel metal1 2574 71 2574 83 7 nResetOut
rlabel metal1 2574 1284 2574 1324 7 Vdd!
rlabel metal1 2574 1260 2574 1272 7 nSDO
rlabel metal1 2574 1233 2574 1245 7 SDI
<< end >>
