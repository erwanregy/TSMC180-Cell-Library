magic
tech tsmc180
timestamp 1701965156
<< nwell >>
rect 0 605 297 1324
<< polysilicon >>
rect 119 703 128 714
rect 119 593 128 605
rect 119 559 128 572
rect 119 494 128 505
<< ndiffusion >>
rect 116 538 119 559
rect 95 505 119 538
rect 128 526 152 559
rect 128 505 131 526
<< pdiffusion >>
rect 115 682 119 703
rect 94 605 119 682
rect 128 626 155 703
rect 128 605 134 626
<< ntransistor >>
rect 119 505 128 559
<< ptransistor >>
rect 119 605 128 703
<< polycontact >>
rect 108 572 129 593
<< ndiffcontact >>
rect 95 538 116 559
rect 131 505 152 526
<< pdiffcontact >>
rect 94 682 115 703
rect 134 605 155 626
<< psubstratetap >>
rect 169 17 204 52
<< nsubstratetap >>
rect 186 1287 221 1322
<< metal1 >>
rect 0 1322 297 1324
rect 0 1305 186 1322
rect 0 1284 94 1305
rect 115 1287 186 1305
rect 221 1287 297 1322
rect 115 1284 297 1287
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 93 703 116 704
rect 93 682 94 703
rect 115 682 116 703
rect 93 681 116 682
rect 134 593 155 605
rect 129 572 155 593
rect 94 559 117 560
rect 94 538 95 559
rect 116 538 117 559
rect 94 537 117 538
rect 240 526 263 527
rect 152 505 241 526
rect 262 505 263 526
rect 240 504 263 505
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 52 241 55
rect 0 17 169 52
rect 204 35 241 52
rect 262 35 297 55
rect 204 17 297 35
rect 0 15 297 17
<< m2contact >>
rect 94 1284 115 1305
rect 94 682 115 703
rect 95 538 116 559
rect 241 505 262 526
rect 241 35 262 55
<< metal2 >>
rect 132 1305 146 1339
rect 132 1284 155 1305
rect 94 703 115 1284
rect 135 608 155 1284
rect 134 559 155 608
rect 116 538 155 559
rect 95 483 116 538
rect 95 462 155 483
rect 135 55 155 462
rect 132 34 155 55
rect 241 55 262 505
rect 132 0 146 34
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal2 132 0 146 0 1 Low
rlabel metal2 132 1339 146 1339 5 Low
<< end >>
