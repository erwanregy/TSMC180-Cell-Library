magic
tech tsmc180
timestamp 1701697717
<< nwell >>
rect 0 605 429 1284
<< polysilicon >>
rect 39 1070 48 1081
rect 110 1070 119 1081
rect 166 1070 175 1081
rect 274 993 283 1079
rect 39 958 48 972
rect 110 958 119 972
rect 166 958 175 972
rect 39 846 48 860
rect 110 846 119 860
rect 166 846 175 860
rect 274 846 283 972
rect 367 768 376 1079
rect 39 703 48 748
rect 110 703 119 748
rect 166 703 175 748
rect 274 703 283 748
rect 367 703 376 747
rect 39 477 48 605
rect 110 477 119 605
rect 166 477 175 605
rect 39 456 76 477
rect 110 456 132 477
rect 166 456 198 477
rect 39 443 48 456
rect 110 443 119 456
rect 166 443 175 456
rect 274 443 283 605
rect 367 443 376 605
rect 39 343 48 389
rect 110 343 119 389
rect 166 343 175 389
rect 274 343 283 388
rect 367 343 376 388
rect 39 275 48 289
rect 110 275 119 289
rect 166 275 175 289
rect 39 207 48 221
rect 110 207 119 221
rect 166 207 175 221
rect 274 207 283 288
rect 39 55 48 153
rect 110 55 119 153
rect 166 55 175 153
rect 274 55 283 186
rect 367 55 376 322
<< ndiffusion >>
rect 36 389 39 443
rect 48 389 110 443
rect 119 389 166 443
rect 175 410 219 443
rect 175 389 198 410
rect 271 421 274 443
rect 250 388 274 421
rect 283 410 318 443
rect 283 389 297 410
rect 283 388 318 389
rect 364 421 367 443
rect 343 388 367 421
rect 376 409 417 443
rect 376 388 396 409
rect 36 289 39 343
rect 48 322 76 343
rect 97 322 110 343
rect 48 289 110 322
rect 119 310 166 343
rect 119 289 132 310
rect 153 289 166 310
rect 175 322 198 343
rect 175 289 219 322
rect 271 322 274 343
rect 250 288 274 322
rect 283 322 297 343
rect 283 288 318 322
rect 36 221 39 275
rect 48 221 110 275
rect 119 242 166 275
rect 119 221 132 242
rect 153 221 166 242
rect 175 221 219 275
rect 36 186 39 207
rect 15 153 39 186
rect 48 175 110 207
rect 48 154 51 175
rect 72 154 110 175
rect 48 153 110 154
rect 119 186 132 207
rect 153 186 166 207
rect 119 153 166 186
rect 175 186 198 207
rect 175 153 219 186
<< pdiffusion >>
rect 15 993 39 1070
rect 36 972 39 993
rect 48 1069 110 1070
rect 48 1048 51 1069
rect 72 1048 110 1069
rect 48 972 110 1048
rect 119 993 166 1070
rect 119 972 132 993
rect 153 972 166 993
rect 175 993 219 1070
rect 175 972 198 993
rect 36 860 39 958
rect 48 860 110 958
rect 119 937 132 958
rect 153 937 166 958
rect 119 860 166 937
rect 175 860 219 958
rect 36 748 39 846
rect 48 769 110 846
rect 48 748 76 769
rect 97 748 110 769
rect 119 825 132 846
rect 153 825 166 846
rect 119 748 166 825
rect 175 769 219 846
rect 175 748 198 769
rect 250 769 274 846
rect 271 748 274 769
rect 283 769 318 846
rect 283 748 297 769
rect 36 605 39 703
rect 48 605 110 703
rect 119 605 166 703
rect 175 682 198 703
rect 175 605 219 682
rect 250 626 274 703
rect 271 605 274 626
rect 283 702 302 703
rect 283 681 297 702
rect 283 605 318 681
rect 343 626 367 703
rect 364 605 367 626
rect 376 682 396 703
rect 376 605 417 682
<< ntransistor >>
rect 39 389 48 443
rect 110 389 119 443
rect 166 389 175 443
rect 274 388 283 443
rect 367 388 376 443
rect 39 289 48 343
rect 110 289 119 343
rect 166 289 175 343
rect 274 288 283 343
rect 39 221 48 275
rect 110 221 119 275
rect 166 221 175 275
rect 39 153 48 207
rect 110 153 119 207
rect 166 153 175 207
<< ptransistor >>
rect 39 972 48 1070
rect 110 972 119 1070
rect 166 972 175 1070
rect 39 860 48 958
rect 110 860 119 958
rect 166 860 175 958
rect 39 748 48 846
rect 110 748 119 846
rect 166 748 175 846
rect 274 748 283 846
rect 39 605 48 703
rect 110 605 119 703
rect 166 605 175 703
rect 274 605 283 703
rect 367 605 376 703
<< polycontact >>
rect 262 972 283 993
rect 355 747 376 768
rect 76 456 97 477
rect 132 456 153 477
rect 198 456 219 477
rect 355 322 376 343
rect 262 186 283 207
<< ndiffcontact >>
rect 15 389 36 443
rect 198 389 219 410
rect 250 421 271 443
rect 297 389 318 410
rect 343 421 364 443
rect 396 388 417 409
rect 15 289 36 343
rect 76 322 97 343
rect 132 289 153 310
rect 198 322 219 343
rect 250 322 271 343
rect 297 322 318 343
rect 15 221 36 275
rect 132 221 153 242
rect 15 186 36 207
rect 51 154 72 175
rect 132 186 153 207
rect 198 186 219 207
<< pdiffcontact >>
rect 15 972 36 993
rect 51 1048 72 1069
rect 132 972 153 993
rect 198 972 219 993
rect 15 860 36 958
rect 132 937 153 958
rect 15 748 36 846
rect 76 748 97 769
rect 132 825 153 846
rect 198 748 219 769
rect 250 748 271 769
rect 297 748 318 769
rect 15 605 36 703
rect 198 682 219 703
rect 250 605 271 626
rect 297 681 318 702
rect 343 605 364 626
rect 396 682 417 703
<< psubstratetap >>
rect 234 18 269 53
<< nsubstratetap >>
rect 235 1285 270 1320
<< metal1 >>
rect 0 1320 429 1324
rect 0 1305 235 1320
rect 0 1284 15 1305
rect 36 1284 51 1305
rect 72 1285 235 1305
rect 270 1285 429 1320
rect 72 1284 429 1285
rect 0 1260 429 1272
rect 0 1233 429 1245
rect 50 1069 73 1070
rect 50 1048 51 1069
rect 72 1048 73 1069
rect 50 1047 73 1048
rect 36 972 132 993
rect 219 972 262 993
rect 14 958 37 959
rect 198 958 219 972
rect 14 860 15 958
rect 36 860 37 958
rect 153 937 219 958
rect 14 859 37 860
rect 14 846 37 847
rect 14 748 15 846
rect 36 825 132 846
rect 36 748 37 825
rect 97 748 198 769
rect 219 748 250 769
rect 318 748 355 768
rect 14 747 37 748
rect 297 747 355 748
rect 297 736 318 747
rect 198 715 318 736
rect 14 703 37 704
rect 14 605 15 703
rect 36 626 37 703
rect 198 703 219 715
rect 395 703 418 704
rect 296 702 319 703
rect 296 681 297 702
rect 318 681 319 702
rect 395 682 396 703
rect 417 682 418 703
rect 395 681 418 682
rect 296 680 319 681
rect 36 605 250 626
rect 271 605 343 626
rect 14 604 37 605
rect 75 477 98 478
rect 75 456 76 477
rect 97 456 98 477
rect 75 455 98 456
rect 131 477 154 478
rect 131 456 132 477
rect 153 456 154 477
rect 131 455 154 456
rect 197 477 220 478
rect 197 456 198 477
rect 219 456 220 477
rect 197 455 220 456
rect 14 443 37 444
rect 14 389 15 443
rect 36 422 250 443
rect 36 389 37 422
rect 271 424 343 443
rect 296 410 319 411
rect 14 388 37 389
rect 198 376 219 389
rect 296 389 297 410
rect 318 389 319 410
rect 296 388 319 389
rect 395 409 418 410
rect 395 388 396 409
rect 417 388 418 409
rect 395 387 418 388
rect 198 355 318 376
rect 14 343 37 344
rect 297 343 318 355
rect 14 289 15 343
rect 36 310 37 343
rect 97 322 198 343
rect 219 322 250 343
rect 318 322 355 343
rect 36 289 132 310
rect 14 288 37 289
rect 14 275 37 276
rect 14 221 15 275
rect 36 221 37 275
rect 153 221 219 242
rect 14 220 37 221
rect 198 207 219 221
rect 36 188 132 207
rect 219 186 262 207
rect 50 175 73 176
rect 50 154 51 175
rect 72 154 73 175
rect 50 153 73 154
rect 0 129 429 141
rect 0 100 429 112
rect 0 71 429 83
rect 0 54 429 55
rect 0 33 15 54
rect 36 33 51 54
rect 72 53 429 54
rect 72 33 234 53
rect 0 18 234 33
rect 269 18 429 53
rect 0 15 429 18
<< m2contact >>
rect 15 1284 36 1305
rect 51 1284 72 1305
rect 51 1048 72 1069
rect 15 860 36 958
rect 15 748 36 846
rect 15 605 36 703
rect 297 681 318 702
rect 396 682 417 703
rect 76 456 97 477
rect 132 456 153 477
rect 198 456 219 477
rect 15 389 36 443
rect 297 389 318 410
rect 396 388 417 409
rect 15 289 36 343
rect 15 221 36 275
rect 51 154 72 175
rect 15 33 36 54
rect 51 33 72 54
<< metal2 >>
rect 99 1324 113 1339
rect 15 958 36 1284
rect 98 1284 113 1324
rect 51 1069 72 1284
rect 92 1033 113 1284
rect 15 846 36 860
rect 15 703 36 748
rect 76 1014 113 1033
rect 132 1081 146 1339
rect 198 1081 212 1339
rect 297 1081 311 1339
rect 396 1081 410 1339
rect 76 477 97 1014
rect 15 343 36 389
rect 15 275 36 289
rect 15 54 36 221
rect 76 210 97 456
rect 132 477 153 1081
rect 76 189 113 210
rect 51 54 72 154
rect 99 0 113 189
rect 132 55 153 456
rect 198 477 219 1081
rect 198 55 219 456
rect 297 702 318 1081
rect 297 410 318 681
rect 297 55 318 389
rect 396 703 417 1081
rect 396 409 417 682
rect 396 55 417 388
rect 132 0 146 55
rect 198 0 212 55
rect 297 0 311 55
rect 396 0 410 55
<< labels >>
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal2 99 1339 113 1339 5 A
rlabel metal2 132 1339 146 1339 5 B
rlabel metal2 198 1339 212 1339 5 Cin
rlabel metal2 297 1339 311 1339 5 Cout
rlabel metal2 396 1339 410 1339 5 S
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 0 15 0 55 3 GND!
rlabel metal2 99 0 113 0 1 A
rlabel metal2 132 0 146 0 1 B
rlabel metal2 198 0 212 0 1 Cin
rlabel metal2 297 0 311 0 1 Cout
rlabel metal2 396 0 410 0 1 S
rlabel metal1 429 1284 429 1324 7 Vdd!
rlabel metal1 429 1260 429 1272 7 ScanReturn
rlabel metal1 429 1233 429 1245 7 Scan
rlabel metal1 429 71 429 83 7 nReset
rlabel metal1 429 100 429 112 7 Clock
rlabel metal1 429 129 429 141 7 Test
rlabel metal1 429 15 429 55 7 GND!
<< end >>
