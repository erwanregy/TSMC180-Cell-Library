magic
tech tsmc180
timestamp 1701965020
<< nwell >>
rect 0 605 429 1324
<< polysilicon >>
rect 39 1071 48 1082
rect 110 1071 119 1082
rect 166 1071 175 1082
rect 274 994 283 1080
rect 39 959 48 973
rect 110 959 119 973
rect 166 959 175 973
rect 39 847 48 861
rect 110 847 119 861
rect 166 847 175 861
rect 274 847 283 973
rect 367 769 376 1080
rect 39 703 48 749
rect 110 703 119 749
rect 166 703 175 749
rect 274 703 283 749
rect 367 703 376 748
rect 39 581 48 605
rect 110 581 119 605
rect 166 581 175 605
rect 39 560 76 581
rect 110 560 132 581
rect 166 560 198 581
rect 39 547 48 560
rect 110 547 119 560
rect 166 547 175 560
rect 274 547 283 605
rect 367 547 376 605
rect 39 447 48 493
rect 110 447 119 493
rect 166 447 175 493
rect 274 447 283 493
rect 367 447 376 493
rect 39 379 48 393
rect 110 379 119 393
rect 166 379 175 393
rect 39 311 48 325
rect 110 311 119 325
rect 166 311 175 325
rect 274 311 283 393
rect 39 55 48 257
rect 110 55 119 257
rect 166 55 175 257
rect 274 55 283 290
rect 367 55 376 426
<< ndiffusion >>
rect 36 493 39 547
rect 48 493 110 547
rect 119 493 166 547
rect 175 514 219 547
rect 175 493 198 514
rect 271 525 274 547
rect 250 493 274 525
rect 283 514 318 547
rect 283 493 297 514
rect 364 525 367 547
rect 343 493 367 525
rect 376 514 417 547
rect 376 493 396 514
rect 36 393 39 447
rect 48 426 76 447
rect 97 426 110 447
rect 48 393 110 426
rect 119 414 166 447
rect 119 393 132 414
rect 153 393 166 414
rect 175 426 198 447
rect 175 393 219 426
rect 271 426 274 447
rect 250 393 274 426
rect 283 426 297 447
rect 283 393 318 426
rect 36 325 39 379
rect 48 325 110 379
rect 119 346 166 379
rect 119 325 132 346
rect 153 325 166 346
rect 175 325 219 379
rect 36 290 39 311
rect 15 257 39 290
rect 48 279 110 311
rect 48 258 51 279
rect 72 258 110 279
rect 48 257 110 258
rect 119 290 132 311
rect 153 290 166 311
rect 119 257 166 290
rect 175 290 198 311
rect 175 257 219 290
<< pdiffusion >>
rect 15 994 39 1071
rect 36 973 39 994
rect 48 1050 51 1071
rect 72 1050 110 1071
rect 48 973 110 1050
rect 119 994 166 1071
rect 119 973 132 994
rect 153 973 166 994
rect 175 994 219 1071
rect 175 973 198 994
rect 36 861 39 959
rect 48 861 110 959
rect 119 938 132 959
rect 153 938 166 959
rect 119 861 166 938
rect 175 861 219 959
rect 36 749 39 847
rect 48 770 110 847
rect 48 749 76 770
rect 97 749 110 770
rect 119 826 132 847
rect 153 826 166 847
rect 119 749 166 826
rect 175 770 219 847
rect 175 749 198 770
rect 250 770 274 847
rect 271 749 274 770
rect 283 770 318 847
rect 283 749 297 770
rect 36 605 39 703
rect 48 605 110 703
rect 119 605 166 703
rect 175 682 198 703
rect 175 605 219 682
rect 250 626 274 703
rect 271 605 274 626
rect 283 682 297 703
rect 283 605 318 682
rect 343 626 367 703
rect 364 605 367 626
rect 376 682 396 703
rect 376 605 417 682
<< ntransistor >>
rect 39 493 48 547
rect 110 493 119 547
rect 166 493 175 547
rect 274 493 283 547
rect 367 493 376 547
rect 39 393 48 447
rect 110 393 119 447
rect 166 393 175 447
rect 274 393 283 447
rect 39 325 48 379
rect 110 325 119 379
rect 166 325 175 379
rect 39 257 48 311
rect 110 257 119 311
rect 166 257 175 311
<< ptransistor >>
rect 39 973 48 1071
rect 110 973 119 1071
rect 166 973 175 1071
rect 39 861 48 959
rect 110 861 119 959
rect 166 861 175 959
rect 39 749 48 847
rect 110 749 119 847
rect 166 749 175 847
rect 274 749 283 847
rect 39 605 48 703
rect 110 605 119 703
rect 166 605 175 703
rect 274 605 283 703
rect 367 605 376 703
<< polycontact >>
rect 262 973 283 994
rect 355 748 376 769
rect 76 560 97 581
rect 132 560 153 581
rect 198 560 219 581
rect 355 426 376 447
rect 262 290 283 311
<< ndiffcontact >>
rect 15 493 36 547
rect 198 493 219 514
rect 250 525 271 547
rect 297 493 318 514
rect 343 525 364 547
rect 396 493 417 514
rect 15 393 36 447
rect 76 426 97 447
rect 132 393 153 414
rect 198 426 219 447
rect 250 426 271 447
rect 297 426 318 447
rect 15 325 36 379
rect 132 325 153 346
rect 15 290 36 311
rect 51 258 72 279
rect 132 290 153 311
rect 198 290 219 311
<< pdiffcontact >>
rect 15 973 36 994
rect 51 1050 72 1071
rect 132 973 153 994
rect 198 973 219 994
rect 15 861 36 959
rect 132 938 153 959
rect 15 749 36 847
rect 76 749 97 770
rect 132 826 153 847
rect 198 749 219 770
rect 250 749 271 770
rect 297 749 318 770
rect 15 605 36 703
rect 198 682 219 703
rect 250 605 271 626
rect 297 682 318 703
rect 343 605 364 626
rect 396 682 417 703
<< psubstratetap >>
rect 234 18 269 53
<< nsubstratetap >>
rect 235 1285 270 1320
<< metal1 >>
rect 0 1320 429 1324
rect 0 1305 235 1320
rect 0 1284 15 1305
rect 36 1284 51 1305
rect 72 1285 235 1305
rect 270 1285 429 1320
rect 72 1284 429 1285
rect 0 1260 429 1272
rect 0 1233 429 1245
rect 50 1071 73 1072
rect 50 1050 51 1071
rect 72 1050 73 1071
rect 50 1049 73 1050
rect 36 973 132 994
rect 219 973 262 994
rect 198 959 219 973
rect 153 938 219 959
rect 36 826 132 847
rect 97 749 198 770
rect 219 749 250 770
rect 318 749 355 769
rect 297 748 355 749
rect 297 737 318 748
rect 198 716 318 737
rect 198 703 219 716
rect 296 703 319 704
rect 296 682 297 703
rect 318 682 319 703
rect 296 681 319 682
rect 395 703 418 704
rect 395 682 396 703
rect 417 682 418 703
rect 395 681 418 682
rect 36 605 250 626
rect 271 605 343 626
rect 75 581 98 582
rect 75 560 76 581
rect 97 560 98 581
rect 75 559 98 560
rect 131 581 154 582
rect 131 560 132 581
rect 153 560 154 581
rect 131 559 154 560
rect 197 581 220 582
rect 197 560 198 581
rect 219 560 220 581
rect 197 559 220 560
rect 36 526 250 547
rect 271 527 343 547
rect 296 514 319 515
rect 198 480 219 493
rect 296 493 297 514
rect 318 493 319 514
rect 296 492 319 493
rect 395 514 418 515
rect 395 493 396 514
rect 417 493 418 514
rect 395 492 418 493
rect 198 459 318 480
rect 297 447 318 459
rect 97 426 198 447
rect 219 426 250 447
rect 318 426 355 447
rect 36 393 132 414
rect 153 325 219 346
rect 198 311 219 325
rect 36 292 132 311
rect 219 290 262 311
rect 50 279 73 280
rect 50 258 51 279
rect 72 258 73 279
rect 50 257 73 258
rect 0 129 429 141
rect 0 100 429 112
rect 0 71 429 83
rect 0 34 15 55
rect 36 34 51 55
rect 72 53 429 55
rect 72 34 234 53
rect 0 18 234 34
rect 269 18 429 53
rect 0 15 429 18
<< m2contact >>
rect 15 1284 36 1305
rect 51 1284 72 1305
rect 51 1050 72 1071
rect 15 861 36 959
rect 15 749 36 847
rect 15 605 36 703
rect 297 682 318 703
rect 396 682 417 703
rect 76 560 97 581
rect 132 560 153 581
rect 198 560 219 581
rect 15 493 36 547
rect 297 493 318 514
rect 396 493 417 514
rect 15 393 36 447
rect 15 325 36 379
rect 51 258 72 279
rect 15 34 36 55
rect 51 34 72 55
<< metal2 >>
rect 99 1324 113 1339
rect 15 959 36 1284
rect 98 1284 113 1324
rect 51 1071 72 1284
rect 92 1036 113 1284
rect 15 847 36 861
rect 15 703 36 749
rect 76 1015 113 1036
rect 132 1082 146 1339
rect 198 1082 212 1339
rect 297 1082 311 1339
rect 396 1082 410 1339
rect 76 581 97 1015
rect 15 447 36 493
rect 15 379 36 393
rect 15 55 36 325
rect 76 314 97 560
rect 132 581 153 1082
rect 76 293 113 314
rect 51 55 72 258
rect 99 0 113 293
rect 132 55 153 560
rect 198 581 219 1082
rect 198 55 219 560
rect 297 703 318 1082
rect 297 514 318 682
rect 297 55 318 493
rect 396 703 417 1082
rect 396 514 417 682
rect 396 55 417 493
rect 132 0 146 55
rect 198 0 212 55
rect 297 0 311 55
rect 396 0 410 55
<< labels >>
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 0 15 0 55 3 GND!
rlabel metal2 99 0 113 0 1 A
rlabel metal2 99 1339 113 1339 5 A
rlabel metal2 132 0 146 0 1 B
rlabel metal2 132 1339 146 1339 5 B
rlabel metal2 198 0 212 0 1 Cin
rlabel metal2 198 1339 212 1339 5 Cin
rlabel metal2 297 0 311 0 1 Cout
rlabel metal2 297 1339 311 1339 5 Cout
rlabel metal2 396 0 410 0 1 S
rlabel metal2 396 1339 410 1339 5 S
rlabel metal1 429 15 429 55 7 GND!
rlabel metal1 429 129 429 141 7 Test
rlabel metal1 429 100 429 112 7 Clock
rlabel metal1 429 71 429 83 7 nReset
rlabel metal1 429 1233 429 1245 7 Scan
rlabel metal1 429 1260 429 1272 7 ScanReturn
rlabel metal1 429 1284 429 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
<< end >>
