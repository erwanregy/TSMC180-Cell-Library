magic
tech tsmc180
timestamp 1701693773
<< nwell >>
rect 0 605 396 1324
<< polysilicon >>
rect 71 927 80 1003
rect 139 927 148 1003
rect 183 927 192 1003
rect 234 927 243 1003
rect 322 927 331 1013
rect 71 722 80 829
rect 71 521 80 624
rect 71 346 80 500
rect 139 388 148 829
rect 71 240 80 292
rect 139 240 148 367
rect 183 612 192 829
rect 183 240 192 591
rect 234 558 243 829
rect 322 798 331 829
rect 329 777 331 798
rect 234 240 243 537
rect 322 273 331 777
rect 322 240 331 252
rect 71 80 80 186
rect 139 118 148 186
rect 183 118 192 186
rect 234 118 243 186
rect 322 150 331 186
<< ndiffusion >>
rect 68 292 71 346
rect 80 292 83 346
rect 68 186 71 240
rect 80 186 114 240
rect 135 186 139 240
rect 148 186 183 240
rect 192 186 207 240
rect 228 186 234 240
rect 243 186 246 240
rect 319 186 322 240
rect 331 186 335 240
<< pdiffusion >>
rect 68 829 71 927
rect 80 829 83 927
rect 104 829 139 927
rect 148 829 156 927
rect 177 829 183 927
rect 192 829 210 927
rect 231 829 234 927
rect 243 829 246 927
rect 319 829 322 927
rect 331 829 335 927
rect 68 624 71 722
rect 80 624 83 722
<< ntransistor >>
rect 71 292 80 346
rect 71 186 80 240
rect 139 186 148 240
rect 183 186 192 240
rect 234 186 243 240
rect 322 186 331 240
<< ptransistor >>
rect 71 829 80 927
rect 139 829 148 927
rect 183 829 192 927
rect 234 829 243 927
rect 322 829 331 927
rect 71 624 80 722
<< polycontact >>
rect 65 500 86 521
rect 127 367 148 388
rect 183 591 204 612
rect 308 777 329 798
rect 228 537 249 558
rect 310 252 331 273
<< ndiffcontact >>
rect 47 292 68 346
rect 83 292 104 346
rect 47 186 68 240
rect 114 186 135 240
rect 207 186 228 240
rect 246 186 267 240
rect 298 186 319 240
rect 335 186 356 240
<< pdiffcontact >>
rect 47 829 68 927
rect 83 829 104 927
rect 156 829 177 927
rect 210 829 231 927
rect 246 829 267 927
rect 298 829 319 927
rect 335 829 356 927
rect 47 624 68 722
rect 83 624 104 722
<< psubstratetap >>
rect 31 30 352 51
<< nsubstratetap >>
rect 42 1293 339 1314
<< metal1 >>
rect 0 1314 396 1324
rect 0 1293 42 1314
rect 339 1293 396 1314
rect 0 1284 396 1293
rect 0 1260 396 1272
rect 0 1233 396 1245
rect 301 987 313 1199
rect 161 975 313 987
rect 161 927 173 975
rect 301 927 313 975
rect 51 793 63 829
rect 86 817 98 829
rect 214 817 226 829
rect 86 805 226 817
rect 249 793 261 829
rect 51 781 308 793
rect 52 752 157 764
rect 52 722 64 752
rect 64 521 87 522
rect 64 500 65 521
rect 86 500 87 521
rect 64 499 87 500
rect 104 388 116 722
rect 182 612 205 613
rect 182 591 183 612
rect 204 591 205 612
rect 182 590 205 591
rect 344 612 356 829
rect 227 558 250 559
rect 227 537 228 558
rect 249 537 250 558
rect 227 536 250 537
rect 104 383 127 388
rect 52 371 127 383
rect 52 346 64 371
rect 104 306 117 325
rect 53 252 159 264
rect 53 240 65 252
rect 147 174 159 252
rect 213 256 310 268
rect 213 240 225 256
rect 344 240 356 593
rect 250 174 262 186
rect 147 162 262 174
rect 0 129 396 141
rect 0 100 396 112
rect 0 71 396 83
rect 0 54 396 55
rect 0 52 300 54
rect 0 51 118 52
rect 137 51 300 52
rect 319 51 396 54
rect 0 30 31 51
rect 352 30 396 51
rect 0 15 396 30
<< m2contact >>
rect 300 1294 319 1313
rect 298 1199 317 1218
rect 156 844 175 863
rect 157 750 176 769
rect 66 501 85 520
rect 184 592 203 611
rect 344 593 363 612
rect 229 538 248 557
rect 117 306 136 325
rect 116 197 135 216
rect 299 195 318 214
rect 118 51 137 52
rect 300 51 319 54
rect 118 33 137 51
rect 300 35 319 51
<< metal2 >>
rect 66 520 80 1339
rect 158 769 172 844
rect 198 611 212 1339
rect 203 592 212 611
rect 66 0 80 501
rect 120 216 134 306
rect 120 52 134 197
rect 198 0 212 592
rect 231 557 245 1339
rect 302 1218 316 1294
rect 231 0 245 538
rect 302 54 316 195
rect 363 0 377 1339
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal2 66 1339 80 1339 5 S
rlabel metal2 66 0 80 0 1 S
rlabel metal2 231 1339 245 1339 5 I1
rlabel metal2 231 0 245 0 1 I1
rlabel metal2 198 0 212 0 1 I0
rlabel metal2 198 1339 212 1339 5 I0
rlabel metal1 396 1233 396 1245 7 Scan
rlabel metal1 396 1260 396 1272 7 ScanReturn
rlabel metal1 396 129 396 141 7 Test
rlabel metal1 396 100 396 112 7 Clock
rlabel metal1 396 71 396 83 7 nReset
rlabel metal2 363 0 377 0 1 Y
rlabel metal2 363 1339 377 1339 5 Y
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal1 396 1284 396 1324 7 Vdd!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 396 15 396 55 7 GND!
<< end >>
