magic
tech tsmc180
timestamp 1701359518
<< nwell >>
rect 546 311 2681 1333
rect 2272 310 2681 311
<< polysilicon >>
rect 1132 966 1141 977
rect 1172 966 1181 977
rect 1212 966 1221 977
rect 1252 966 1261 977
rect 937 620 946 631
rect 977 620 986 631
rect 1017 620 1026 631
rect 1057 620 1066 631
rect 823 568 832 580
rect 861 568 870 580
rect 750 529 759 543
rect 613 515 622 529
rect 613 358 622 417
rect 750 359 759 417
rect 823 359 832 417
rect 613 284 622 337
rect 750 284 759 338
rect 823 303 832 338
rect 861 303 870 417
rect 937 357 946 416
rect 823 294 870 303
rect 823 284 832 294
rect 861 284 870 294
rect 937 306 946 336
rect 977 306 986 416
rect 1017 306 1026 416
rect 1057 306 1066 416
rect 1786 964 1795 975
rect 1826 964 1835 975
rect 1866 964 1875 975
rect 1906 964 1915 975
rect 1591 618 1600 629
rect 1631 618 1640 629
rect 1671 618 1680 629
rect 1711 618 1720 629
rect 1477 566 1486 578
rect 1515 566 1524 578
rect 1404 527 1413 541
rect 1132 356 1141 415
rect 937 297 1066 306
rect 937 284 946 297
rect 977 284 986 297
rect 1017 284 1026 297
rect 1057 284 1066 297
rect 1132 313 1141 335
rect 1172 313 1181 415
rect 1212 313 1221 415
rect 1252 313 1261 415
rect 1404 359 1413 415
rect 1477 359 1486 415
rect 1132 304 1261 313
rect 1132 284 1141 304
rect 1172 284 1181 304
rect 1212 284 1221 304
rect 1252 284 1261 304
rect 1404 284 1413 338
rect 1477 303 1486 338
rect 1515 303 1524 415
rect 1591 357 1600 414
rect 1477 294 1524 303
rect 1477 284 1486 294
rect 1515 284 1524 294
rect 1591 306 1600 336
rect 1631 306 1640 414
rect 1671 306 1680 414
rect 1711 306 1720 414
rect 2435 962 2444 973
rect 2475 962 2484 973
rect 2515 962 2524 973
rect 2555 962 2564 973
rect 2240 616 2249 627
rect 2280 616 2289 627
rect 2320 616 2329 627
rect 2360 616 2369 627
rect 2126 564 2135 576
rect 2164 564 2173 576
rect 2053 525 2062 539
rect 1786 356 1795 413
rect 1591 297 1720 306
rect 1591 284 1600 297
rect 1631 284 1640 297
rect 1671 284 1680 297
rect 1711 284 1720 297
rect 1786 313 1795 335
rect 1826 313 1835 413
rect 1866 313 1875 413
rect 1906 313 1915 413
rect 2053 359 2062 413
rect 2126 359 2135 413
rect 1786 304 1915 313
rect 1786 284 1795 304
rect 1826 284 1835 304
rect 1866 284 1875 304
rect 1906 284 1915 304
rect 2053 284 2062 338
rect 2126 303 2135 338
rect 2164 303 2173 413
rect 2240 357 2249 412
rect 2126 294 2173 303
rect 2126 284 2135 294
rect 2164 284 2173 294
rect 2240 306 2249 336
rect 2280 306 2289 412
rect 2320 306 2329 412
rect 2360 306 2369 412
rect 2435 356 2444 411
rect 2240 297 2369 306
rect 2240 284 2249 297
rect 2280 284 2289 297
rect 2320 284 2329 297
rect 2360 284 2369 297
rect 2435 313 2444 335
rect 2475 313 2484 411
rect 2515 313 2524 411
rect 2555 313 2564 411
rect 2435 304 2564 313
rect 2435 284 2444 304
rect 2475 284 2484 304
rect 2515 284 2524 304
rect 2555 284 2564 304
rect 750 231 759 242
rect 613 219 622 230
rect 823 217 832 228
rect 861 217 870 228
rect 937 197 946 208
rect 977 197 986 208
rect 1017 197 1026 208
rect 1057 197 1066 208
rect 1404 231 1413 242
rect 1477 217 1486 228
rect 1515 217 1524 228
rect 1591 197 1600 208
rect 1631 197 1640 208
rect 1671 197 1680 208
rect 1711 197 1720 208
rect 2053 231 2062 242
rect 2126 217 2135 228
rect 2164 217 2173 228
rect 2240 197 2249 208
rect 2280 197 2289 208
rect 2320 197 2329 208
rect 2360 197 2369 208
rect 1132 65 1141 77
rect 1172 65 1181 77
rect 1212 65 1221 77
rect 1252 65 1261 77
rect 1786 65 1795 77
rect 1826 65 1835 77
rect 1866 65 1875 77
rect 1906 65 1915 77
rect 2435 65 2444 77
rect 2475 65 2484 77
rect 2515 65 2524 77
rect 2555 65 2564 77
<< ndiffusion >>
rect 608 230 613 284
rect 622 230 627 284
rect 745 242 750 284
rect 759 242 764 284
rect 820 228 823 284
rect 832 228 836 284
rect 857 228 861 284
rect 870 228 875 284
rect 932 208 937 284
rect 946 208 951 284
rect 972 208 977 284
rect 986 208 991 284
rect 1012 208 1017 284
rect 1026 208 1031 284
rect 1052 208 1057 284
rect 1066 208 1071 284
rect 1127 77 1132 284
rect 1141 77 1146 284
rect 1167 77 1172 284
rect 1181 77 1186 284
rect 1207 77 1212 284
rect 1221 77 1226 284
rect 1247 77 1252 284
rect 1261 77 1266 284
rect 1399 242 1404 284
rect 1413 242 1418 284
rect 1474 228 1477 284
rect 1486 228 1490 284
rect 1511 228 1515 284
rect 1524 228 1529 284
rect 1586 208 1591 284
rect 1600 208 1605 284
rect 1626 208 1631 284
rect 1640 208 1645 284
rect 1666 208 1671 284
rect 1680 208 1685 284
rect 1706 208 1711 284
rect 1720 208 1725 284
rect 1781 77 1786 284
rect 1795 77 1800 284
rect 1821 77 1826 284
rect 1835 77 1840 284
rect 1861 77 1866 284
rect 1875 77 1880 284
rect 1901 77 1906 284
rect 1915 77 1920 284
rect 2048 242 2053 284
rect 2062 242 2067 284
rect 2123 228 2126 284
rect 2135 228 2139 284
rect 2160 228 2164 284
rect 2173 228 2178 284
rect 2235 208 2240 284
rect 2249 208 2254 284
rect 2275 208 2280 284
rect 2289 208 2294 284
rect 2315 208 2320 284
rect 2329 208 2334 284
rect 2355 208 2360 284
rect 2369 208 2374 284
rect 2430 77 2435 284
rect 2444 77 2449 284
rect 2470 77 2475 284
rect 2484 77 2489 284
rect 2510 77 2515 284
rect 2524 77 2529 284
rect 2550 77 2555 284
rect 2564 77 2569 284
<< pdiffusion >>
rect 608 417 613 515
rect 622 417 627 515
rect 745 417 750 529
rect 759 417 764 529
rect 820 417 823 568
rect 832 417 836 568
rect 857 417 861 568
rect 870 417 876 568
rect 932 416 937 620
rect 946 416 951 620
rect 972 416 977 620
rect 986 416 991 620
rect 1012 416 1017 620
rect 1026 416 1031 620
rect 1052 416 1057 620
rect 1066 416 1071 620
rect 1127 415 1132 966
rect 1141 415 1146 966
rect 1167 415 1172 966
rect 1181 415 1186 966
rect 1207 415 1212 966
rect 1221 415 1226 966
rect 1247 415 1252 966
rect 1261 415 1266 966
rect 1399 415 1404 527
rect 1413 415 1418 527
rect 1474 415 1477 566
rect 1486 415 1490 566
rect 1511 415 1515 566
rect 1524 415 1530 566
rect 1586 414 1591 618
rect 1600 414 1605 618
rect 1626 414 1631 618
rect 1640 414 1645 618
rect 1666 414 1671 618
rect 1680 414 1685 618
rect 1706 414 1711 618
rect 1720 414 1725 618
rect 1781 413 1786 964
rect 1795 413 1800 964
rect 1821 413 1826 964
rect 1835 413 1840 964
rect 1861 413 1866 964
rect 1875 413 1880 964
rect 1901 413 1906 964
rect 1915 413 1920 964
rect 2048 413 2053 525
rect 2062 413 2067 525
rect 2123 413 2126 564
rect 2135 413 2139 564
rect 2160 413 2164 564
rect 2173 413 2179 564
rect 2235 412 2240 616
rect 2249 412 2254 616
rect 2275 412 2280 616
rect 2289 412 2294 616
rect 2315 412 2320 616
rect 2329 412 2334 616
rect 2355 412 2360 616
rect 2369 412 2374 616
rect 2430 411 2435 962
rect 2444 411 2449 962
rect 2470 411 2475 962
rect 2484 411 2489 962
rect 2510 411 2515 962
rect 2524 411 2529 962
rect 2550 411 2555 962
rect 2564 411 2569 962
<< ntransistor >>
rect 613 230 622 284
rect 750 242 759 284
rect 823 228 832 284
rect 861 228 870 284
rect 937 208 946 284
rect 977 208 986 284
rect 1017 208 1026 284
rect 1057 208 1066 284
rect 1132 77 1141 284
rect 1172 77 1181 284
rect 1212 77 1221 284
rect 1252 77 1261 284
rect 1404 242 1413 284
rect 1477 228 1486 284
rect 1515 228 1524 284
rect 1591 208 1600 284
rect 1631 208 1640 284
rect 1671 208 1680 284
rect 1711 208 1720 284
rect 1786 77 1795 284
rect 1826 77 1835 284
rect 1866 77 1875 284
rect 1906 77 1915 284
rect 2053 242 2062 284
rect 2126 228 2135 284
rect 2164 228 2173 284
rect 2240 208 2249 284
rect 2280 208 2289 284
rect 2320 208 2329 284
rect 2360 208 2369 284
rect 2435 77 2444 284
rect 2475 77 2484 284
rect 2515 77 2524 284
rect 2555 77 2564 284
<< ptransistor >>
rect 613 417 622 515
rect 750 417 759 529
rect 823 417 832 568
rect 861 417 870 568
rect 937 416 946 620
rect 977 416 986 620
rect 1017 416 1026 620
rect 1057 416 1066 620
rect 1132 415 1141 966
rect 1172 415 1181 966
rect 1212 415 1221 966
rect 1252 415 1261 966
rect 1404 415 1413 527
rect 1477 415 1486 566
rect 1515 415 1524 566
rect 1591 414 1600 618
rect 1631 414 1640 618
rect 1671 414 1680 618
rect 1711 414 1720 618
rect 1786 413 1795 964
rect 1826 413 1835 964
rect 1866 413 1875 964
rect 1906 413 1915 964
rect 2053 413 2062 525
rect 2126 413 2135 564
rect 2164 413 2173 564
rect 2240 412 2249 616
rect 2280 412 2289 616
rect 2320 412 2329 616
rect 2360 412 2369 616
rect 2435 411 2444 962
rect 2475 411 2484 962
rect 2515 411 2524 962
rect 2555 411 2564 962
<< polycontact >>
rect 613 337 634 358
rect 738 338 759 359
rect 810 338 832 359
rect 925 336 946 357
rect 1120 335 1141 356
rect 1392 338 1413 359
rect 1464 338 1486 359
rect 1579 336 1600 357
rect 1774 335 1795 356
rect 2041 338 2062 359
rect 2113 338 2135 359
rect 2228 336 2249 357
rect 2423 335 2444 356
<< ndiffcontact >>
rect 587 230 608 284
rect 627 230 648 284
rect 724 242 745 284
rect 764 242 785 284
rect 799 228 820 284
rect 836 228 857 284
rect 875 228 896 284
rect 911 208 932 284
rect 951 208 972 284
rect 991 208 1012 284
rect 1031 208 1052 284
rect 1071 208 1092 284
rect 1106 77 1127 284
rect 1146 77 1167 284
rect 1186 77 1207 284
rect 1226 77 1247 284
rect 1266 77 1287 284
rect 1378 242 1399 284
rect 1418 242 1439 284
rect 1453 228 1474 284
rect 1490 228 1511 284
rect 1529 228 1550 284
rect 1565 208 1586 284
rect 1605 208 1626 284
rect 1645 208 1666 284
rect 1685 208 1706 284
rect 1725 208 1746 284
rect 1760 77 1781 284
rect 1800 77 1821 284
rect 1840 77 1861 284
rect 1880 77 1901 284
rect 1920 77 1941 284
rect 2027 242 2048 284
rect 2067 242 2088 284
rect 2102 228 2123 284
rect 2139 228 2160 284
rect 2178 228 2199 284
rect 2214 208 2235 284
rect 2254 208 2275 284
rect 2294 208 2315 284
rect 2334 208 2355 284
rect 2374 208 2395 284
rect 2409 77 2430 284
rect 2449 77 2470 284
rect 2489 77 2510 284
rect 2529 77 2550 284
rect 2569 77 2590 284
<< pdiffcontact >>
rect 587 417 608 515
rect 627 417 648 515
rect 724 417 745 529
rect 764 417 785 529
rect 799 417 820 568
rect 836 417 857 568
rect 876 417 897 568
rect 911 416 932 620
rect 951 416 972 620
rect 991 416 1012 620
rect 1031 416 1052 620
rect 1071 416 1092 620
rect 1106 415 1127 966
rect 1146 415 1167 966
rect 1186 415 1207 966
rect 1226 415 1247 966
rect 1266 415 1287 966
rect 1378 415 1399 527
rect 1418 415 1439 527
rect 1453 415 1474 566
rect 1490 415 1511 566
rect 1530 415 1551 566
rect 1565 414 1586 618
rect 1605 414 1626 618
rect 1645 414 1666 618
rect 1685 414 1706 618
rect 1725 414 1746 618
rect 1760 413 1781 964
rect 1800 413 1821 964
rect 1840 413 1861 964
rect 1880 413 1901 964
rect 1920 413 1941 964
rect 2027 413 2048 525
rect 2067 413 2088 525
rect 2102 413 2123 564
rect 2139 413 2160 564
rect 2179 413 2200 564
rect 2214 412 2235 616
rect 2254 412 2275 616
rect 2294 412 2315 616
rect 2334 412 2355 616
rect 2374 412 2395 616
rect 2409 411 2430 962
rect 2449 411 2470 962
rect 2489 411 2510 962
rect 2529 411 2550 962
rect 2569 411 2590 962
<< psubstratetap >>
rect 810 18 845 53
rect 876 19 911 54
rect 987 16 1022 51
rect 1177 15 1212 50
rect 1342 15 1377 50
rect 1412 15 1447 50
rect 1625 16 1660 51
rect 1734 15 1769 50
rect 1927 15 1962 50
rect 2191 15 2226 50
rect 2354 16 2389 51
rect 2482 15 2517 50
rect 2556 15 2591 50
rect 2612 15 2647 50
<< nsubstratetap >>
rect 657 1284 692 1319
rect 832 1289 867 1324
rect 1136 1287 1171 1322
rect 1406 1286 1441 1321
rect 1593 1288 1628 1323
rect 1784 1284 1819 1319
rect 1878 1289 1913 1324
rect 2127 1286 2162 1321
rect 2247 1287 2282 1322
rect 2325 1289 2360 1324
rect 2519 1288 2554 1323
rect 2609 1286 2644 1321
<< metal1 >>
rect 219 1319 832 1324
rect 219 1313 657 1319
rect 219 1292 627 1313
rect 648 1292 657 1313
rect 219 1284 657 1292
rect 692 1314 832 1319
rect 692 1313 799 1314
rect 692 1292 724 1313
rect 745 1293 799 1313
rect 820 1293 832 1314
rect 745 1292 832 1293
rect 692 1289 832 1292
rect 867 1323 1878 1324
rect 867 1322 1593 1323
rect 867 1317 1136 1322
rect 867 1296 876 1317
rect 897 1313 1136 1317
rect 897 1312 991 1313
rect 897 1296 911 1312
rect 867 1291 911 1296
rect 932 1292 991 1312
rect 1012 1292 1071 1313
rect 1092 1292 1106 1313
rect 1127 1292 1136 1313
rect 932 1291 1136 1292
rect 867 1289 1136 1291
rect 692 1287 1136 1289
rect 1171 1321 1593 1322
rect 1171 1315 1406 1321
rect 1171 1313 1378 1315
rect 1171 1292 1186 1313
rect 1207 1292 1266 1313
rect 1287 1296 1378 1313
rect 1399 1296 1406 1315
rect 1287 1292 1406 1296
rect 1171 1287 1406 1292
rect 692 1286 1406 1287
rect 1441 1313 1593 1321
rect 1441 1309 1565 1313
rect 1441 1290 1453 1309
rect 1474 1290 1530 1309
rect 1551 1294 1565 1309
rect 1586 1294 1593 1313
rect 1551 1290 1593 1294
rect 1441 1288 1593 1290
rect 1628 1319 1878 1323
rect 1628 1314 1784 1319
rect 1628 1313 1760 1314
rect 1628 1310 1725 1313
rect 1628 1291 1645 1310
rect 1666 1294 1725 1310
rect 1746 1295 1760 1313
rect 1781 1295 1784 1314
rect 1746 1294 1784 1295
rect 1666 1291 1784 1294
rect 1628 1288 1784 1291
rect 1441 1286 1784 1288
rect 692 1284 1784 1286
rect 1819 1313 1878 1319
rect 1819 1294 1840 1313
rect 1861 1294 1878 1313
rect 1819 1289 1878 1294
rect 1913 1322 2325 1324
rect 1913 1321 2247 1322
rect 1913 1314 2127 1321
rect 1913 1295 1920 1314
rect 1941 1295 2027 1314
rect 2048 1313 2127 1314
rect 2048 1295 2102 1313
rect 1913 1294 2102 1295
rect 2123 1294 2127 1313
rect 1913 1289 2127 1294
rect 1819 1286 2127 1289
rect 2162 1314 2247 1321
rect 2162 1312 2214 1314
rect 2162 1293 2179 1312
rect 2200 1295 2214 1312
rect 2235 1295 2247 1314
rect 2200 1293 2247 1295
rect 2162 1287 2247 1293
rect 2282 1308 2325 1322
rect 2282 1289 2294 1308
rect 2315 1289 2325 1308
rect 2360 1314 2519 1324
rect 2360 1295 2374 1314
rect 2395 1295 2409 1314
rect 2430 1311 2519 1314
rect 2430 1295 2489 1311
rect 2360 1292 2489 1295
rect 2510 1292 2519 1311
rect 2360 1289 2519 1292
rect 2282 1288 2519 1289
rect 2554 1321 2699 1324
rect 2554 1316 2609 1321
rect 2554 1297 2569 1316
rect 2590 1297 2609 1316
rect 2554 1288 2609 1297
rect 2282 1287 2609 1288
rect 2162 1286 2609 1287
rect 2644 1286 2699 1321
rect 1819 1284 2699 1286
rect 446 1257 557 1269
rect 682 1260 2699 1272
rect 2620 1237 2699 1245
rect 447 1233 2699 1237
rect 447 1225 2632 1233
rect 479 1190 691 1202
rect 512 1156 1345 1168
rect 545 1130 1994 1142
rect 1320 1096 2663 1108
rect 1980 1054 2638 1066
rect 1106 966 1127 986
rect 1186 966 1207 986
rect 1266 966 1287 986
rect 627 515 648 568
rect 724 529 745 712
rect 799 568 820 712
rect 876 568 897 711
rect 911 620 932 711
rect 991 620 1012 711
rect 1071 620 1092 711
rect 587 355 601 417
rect 575 340 601 355
rect 587 284 601 340
rect 634 341 659 353
rect 714 342 738 354
rect 771 356 785 417
rect 771 341 810 356
rect 771 284 785 341
rect 845 352 857 417
rect 956 404 969 416
rect 1036 404 1048 416
rect 1760 964 1781 984
rect 1840 964 1861 984
rect 1920 964 1941 984
rect 1378 527 1399 710
rect 1453 566 1474 710
rect 1530 566 1551 709
rect 1565 618 1586 709
rect 1645 618 1666 709
rect 1725 618 1746 709
rect 956 391 1048 404
rect 845 340 925 352
rect 845 284 857 340
rect 1035 351 1048 391
rect 1151 403 1164 415
rect 1231 403 1243 415
rect 1151 390 1282 403
rect 1267 356 1282 390
rect 1035 339 1120 351
rect 1035 309 1048 339
rect 1267 341 1301 356
rect 1267 323 1282 341
rect 1368 342 1392 354
rect 1425 356 1439 415
rect 1425 341 1464 356
rect 958 296 1048 309
rect 958 284 971 296
rect 1035 284 1048 296
rect 1153 310 1282 323
rect 1153 284 1166 310
rect 1230 284 1243 310
rect 1425 284 1439 341
rect 1499 352 1511 415
rect 1610 402 1623 414
rect 1690 402 1702 414
rect 2409 962 2430 982
rect 2489 962 2510 982
rect 2569 962 2590 982
rect 2027 525 2048 708
rect 2102 564 2123 708
rect 2179 564 2200 707
rect 2214 616 2235 707
rect 2294 616 2315 707
rect 2374 616 2395 707
rect 1610 389 1702 402
rect 1499 340 1579 352
rect 1499 284 1511 340
rect 1689 351 1702 389
rect 1805 401 1818 413
rect 1885 401 1897 413
rect 1805 388 1936 401
rect 1689 339 1774 351
rect 1689 309 1702 339
rect 1921 348 1936 388
rect 1921 333 1959 348
rect 1921 323 1936 333
rect 2017 342 2041 354
rect 2074 356 2088 413
rect 2074 341 2113 356
rect 1612 296 1702 309
rect 1612 284 1625 296
rect 1689 284 1702 296
rect 1807 310 1936 323
rect 1807 284 1820 310
rect 1884 284 1897 310
rect 2074 284 2088 341
rect 2148 352 2160 413
rect 2259 400 2272 412
rect 2339 400 2351 412
rect 2259 387 2351 400
rect 2148 340 2228 352
rect 2148 284 2160 340
rect 2338 351 2351 387
rect 2454 399 2467 411
rect 2534 399 2546 411
rect 2454 386 2585 399
rect 2338 339 2423 351
rect 2338 309 2351 339
rect 2570 323 2585 386
rect 2261 296 2351 309
rect 2261 284 2274 296
rect 2338 284 2351 296
rect 2456 322 2585 323
rect 2456 310 2614 322
rect 2456 284 2469 310
rect 2533 284 2546 310
rect 627 219 648 230
rect 626 55 647 219
rect 724 55 745 242
rect 799 55 820 228
rect 875 55 896 228
rect 913 55 930 208
rect 991 55 1012 208
rect 1072 55 1089 208
rect 1108 55 1123 77
rect 1189 55 1204 77
rect 1267 76 1283 77
rect 1268 55 1283 76
rect 1378 55 1399 242
rect 1453 55 1474 228
rect 1529 55 1550 228
rect 1567 55 1584 208
rect 1645 55 1666 208
rect 1726 55 1743 208
rect 1762 55 1777 77
rect 1843 55 1858 77
rect 1921 76 1937 77
rect 1922 55 1937 76
rect 2027 55 2048 242
rect 2102 55 2123 228
rect 2178 55 2199 228
rect 2216 55 2233 208
rect 2294 55 2315 208
rect 2375 55 2392 208
rect 2602 83 2614 310
rect 2626 112 2638 1054
rect 2651 141 2663 1096
rect 2651 129 2699 141
rect 2626 100 2699 112
rect 2411 55 2426 77
rect 2492 55 2507 77
rect 2570 76 2586 77
rect 2571 55 2586 76
rect 2602 71 2699 83
rect 626 54 2699 55
rect 626 53 876 54
rect 626 18 810 53
rect 845 19 876 53
rect 911 51 2699 54
rect 911 19 987 51
rect 845 18 987 19
rect 626 16 987 18
rect 1022 50 1625 51
rect 1022 16 1177 50
rect 626 15 1177 16
rect 1212 15 1342 50
rect 1377 15 1412 50
rect 1447 16 1625 50
rect 1660 50 2354 51
rect 1660 16 1734 50
rect 1447 15 1734 16
rect 1769 15 1927 50
rect 1962 15 2191 50
rect 2226 16 2354 50
rect 2389 50 2699 51
rect 2389 16 2482 50
rect 2226 15 2482 16
rect 2517 15 2556 50
rect 2591 15 2612 50
rect 2647 15 2699 50
<< m2contact >>
rect 179 1284 219 1324
rect 627 1292 648 1313
rect 724 1292 745 1313
rect 799 1293 820 1314
rect 876 1296 897 1317
rect 911 1291 932 1312
rect 991 1292 1012 1313
rect 1071 1292 1092 1313
rect 1106 1292 1127 1313
rect 1186 1292 1207 1313
rect 1266 1292 1287 1313
rect 1378 1296 1399 1315
rect 1453 1290 1474 1309
rect 1530 1290 1551 1309
rect 1565 1294 1586 1313
rect 1645 1291 1666 1310
rect 1725 1294 1746 1313
rect 1760 1295 1781 1314
rect 1840 1294 1861 1313
rect 1920 1295 1941 1314
rect 2027 1295 2048 1314
rect 2102 1294 2123 1313
rect 2179 1293 2200 1312
rect 2214 1295 2235 1314
rect 2294 1289 2315 1308
rect 2374 1295 2395 1314
rect 2409 1295 2430 1314
rect 2489 1292 2510 1311
rect 2569 1297 2590 1316
rect 427 1253 446 1272
rect 557 1253 576 1272
rect 663 1253 682 1272
rect 428 1218 447 1237
rect 460 1185 479 1204
rect 691 1187 710 1206
rect 493 1152 512 1171
rect 1345 1155 1364 1174
rect 526 1123 545 1142
rect 1994 1127 2013 1146
rect 1301 1090 1320 1109
rect 1961 1054 1980 1073
rect 1106 986 1127 1007
rect 1186 986 1207 1007
rect 1266 986 1287 1007
rect 724 712 745 733
rect 627 568 648 589
rect 799 712 820 733
rect 876 711 897 732
rect 911 711 932 732
rect 991 711 1012 732
rect 1071 711 1092 732
rect 556 338 575 357
rect 659 338 678 357
rect 695 339 714 358
rect 1760 984 1781 1005
rect 1840 984 1861 1005
rect 1920 984 1941 1005
rect 1378 710 1399 731
rect 1453 710 1474 731
rect 1530 709 1551 730
rect 1565 709 1586 730
rect 1645 709 1666 730
rect 1725 709 1746 730
rect 1301 338 1320 357
rect 1349 339 1368 358
rect 2409 982 2430 1003
rect 2489 982 2510 1003
rect 2569 982 2590 1003
rect 2027 708 2048 729
rect 2102 708 2123 729
rect 2179 707 2200 728
rect 2214 707 2235 728
rect 2294 707 2315 728
rect 2374 707 2395 728
rect 1959 331 1978 350
rect 1998 339 2017 358
<< metal2 >>
rect 0 1324 400 1339
rect 0 1284 179 1324
rect 219 1284 400 1324
rect 0 0 400 1284
rect 429 1272 443 1339
rect 429 0 443 1218
rect 462 1204 476 1339
rect 462 0 476 1185
rect 495 1171 509 1339
rect 495 0 509 1152
rect 528 1142 542 1339
rect 528 0 542 1123
rect 559 357 573 1253
rect 627 589 648 1292
rect 663 357 677 1253
rect 696 358 710 1187
rect 724 733 745 1292
rect 799 733 820 1293
rect 876 732 897 1296
rect 911 732 932 1291
rect 991 732 1012 1292
rect 1071 732 1092 1292
rect 1106 1007 1127 1292
rect 1186 1007 1207 1292
rect 1266 1007 1287 1292
rect 1301 357 1315 1090
rect 1350 358 1364 1155
rect 1378 731 1399 1296
rect 1453 731 1474 1290
rect 1530 730 1551 1290
rect 1565 730 1586 1294
rect 1645 730 1666 1291
rect 1725 730 1746 1294
rect 1760 1005 1781 1295
rect 1840 1005 1861 1294
rect 1920 1005 1941 1295
rect 1962 752 1978 1054
rect 1964 350 1978 752
rect 1999 358 2013 1127
rect 2027 729 2048 1295
rect 2102 729 2123 1294
rect 2179 728 2200 1293
rect 2214 728 2235 1295
rect 2294 728 2315 1289
rect 2374 728 2395 1295
rect 2409 1003 2430 1295
rect 2489 1003 2510 1292
rect 2569 1003 2590 1297
<< labels >>
rlabel metal2 0 0 400 0 1 Vdd!
rlabel metal2 462 0 476 0 1 Test
rlabel metal2 495 0 509 0 1 Clock
rlabel metal2 528 0 542 0 1 nReset
rlabel metal2 429 0 443 0 1 SDI
rlabel metal2 0 1339 400 1339 5 Vdd!
rlabel metal2 429 1339 443 1339 5 SDO
rlabel metal2 495 1339 509 1339 5 Clock
rlabel metal2 462 1339 476 1339 5 Test
rlabel metal2 528 1339 542 1339 5 nReset
rlabel metal1 2699 15 2699 55 7 GND!
rlabel metal1 2699 129 2699 141 7 TestOut
rlabel metal1 2699 100 2699 112 7 ClockOut
rlabel metal1 2699 71 2699 83 7 nResetOut
rlabel metal1 2699 1284 2699 1324 7 Vdd!
rlabel metal1 2699 1260 2699 1272 7 nSDO
rlabel metal1 2699 1233 2699 1245 7 SDI
<< end >>
