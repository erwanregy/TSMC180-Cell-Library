magic
tech tsmc180
timestamp 1701692953
<< nwell >>
rect 0 605 297 1284
<< polysilicon >>
rect 119 706 128 717
rect 119 596 128 607
rect 119 562 128 575
rect 119 497 128 508
<< ndiffusion >>
rect 116 541 119 562
rect 95 508 119 541
rect 128 529 152 562
rect 128 508 131 529
<< pdiffusion >>
rect 115 685 119 706
rect 94 607 119 685
rect 128 628 155 706
rect 128 607 134 628
<< ntransistor >>
rect 119 508 128 562
<< ptransistor >>
rect 119 607 128 706
<< polycontact >>
rect 108 575 129 596
<< ndiffcontact >>
rect 95 541 116 562
rect 131 508 152 529
<< pdiffcontact >>
rect 94 685 115 706
rect 134 607 155 628
<< psubstratetap >>
rect 169 17 204 52
<< nsubstratetap >>
rect 186 1287 221 1322
<< metal1 >>
rect 0 1322 297 1324
rect 0 1306 186 1322
rect 0 1285 94 1306
rect 115 1287 186 1306
rect 221 1287 297 1322
rect 115 1285 297 1287
rect 0 1284 297 1285
rect 0 1260 297 1272
rect 0 1233 297 1245
rect 93 706 116 707
rect 93 685 94 706
rect 115 685 116 706
rect 93 684 116 685
rect 134 596 155 607
rect 129 575 155 596
rect 94 562 117 563
rect 94 541 95 562
rect 116 541 117 562
rect 94 540 117 541
rect 240 529 263 530
rect 152 508 241 529
rect 262 508 263 529
rect 240 507 263 508
rect 0 129 297 141
rect 0 100 297 112
rect 0 71 297 83
rect 0 54 297 55
rect 0 52 241 54
rect 0 17 169 52
rect 204 34 241 52
rect 262 34 297 54
rect 204 17 297 34
rect 0 15 297 17
<< m2contact >>
rect 94 1285 115 1306
rect 94 685 115 706
rect 95 541 116 562
rect 241 508 262 529
rect 241 34 262 54
<< metal2 >>
rect 94 706 115 1285
rect 132 1305 146 1339
rect 132 1284 155 1305
rect 135 610 155 1284
rect 134 562 155 610
rect 116 541 155 562
rect 95 486 116 541
rect 95 465 155 486
rect 135 55 155 465
rect 132 34 155 55
rect 241 54 262 508
rect 132 0 146 34
<< labels >>
rlabel metal1 0 1260 0 1272 3 ScanReturn
rlabel metal1 0 1233 0 1245 3 Scan
rlabel metal1 297 1260 297 1272 7 ScanReturn
rlabel metal1 297 1233 297 1245 7 Scan
rlabel metal1 297 129 297 141 7 Test
rlabel metal1 297 100 297 112 7 Clock
rlabel metal1 297 71 297 83 7 nReset
rlabel metal1 297 15 297 55 7 GND!
rlabel metal1 0 15 0 55 3 GND!
rlabel metal1 0 71 0 83 3 nReset
rlabel metal1 0 100 0 112 3 Clock
rlabel metal1 0 129 0 141 3 Test
rlabel metal1 297 1284 297 1324 7 Vdd!
rlabel metal1 0 1284 0 1324 3 Vdd!
rlabel metal2 132 0 146 0 1 High
rlabel metal2 132 1339 146 1339 5 High
<< end >>